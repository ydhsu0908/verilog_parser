
module HS_TXCTL ( DATA_TX, TXVALID, TXREADY, CLK60M, TXSTART, STSRST_, TX_PID, 
    CRC, TXSOF, TOKEN, DATPKT, HANDSHK, SPLIT, TRST_, DIS_STUFF, MAXLEN, 
    HOSTDAT, TXCRCEN, TXCRCRST, ADRENDPS, USBPOP, PKTXEND, TXCRCDAT, TXBCNT, 
    TEST_J, TEST_K, TEST_PACKET, TEST_EYE, TXCRCPHASE, SL_TXDATASEL, 
    SL_TXFIXDATA, SL_FORCE_CRC, SL_FORCE_STUFF, SOF_DISCONN_CHK, 
    DIS_NARROW_SOF, SOF_DISCONN, TURN_PARM, FORCE_CRCERR, EN_UTM_SPDUP, 
    TURNCNT_EN, ATPG_ENI );
output [7:0] DATA_TX;
input  [7:0] TX_PID;
input  [7:0] HOSTDAT;
input  [18:0] ADRENDPS;
input  [2:0] SL_TXDATASEL;
input  [3:0] TURN_PARM;
input  [15:0] CRC;
output [7:0] TXCRCDAT;
input  [10:0] MAXLEN;
input  [7:0] SL_TXFIXDATA;
output [10:0] TXBCNT;
input  TXREADY, CLK60M, TXSTART, STSRST_, TXSOF, TOKEN, DATPKT, HANDSHK, SPLIT, 
    TRST_, TEST_J, TEST_K, TEST_PACKET, TEST_EYE, SL_FORCE_CRC, SL_FORCE_STUFF, 
    SOF_DISCONN_CHK, DIS_NARROW_SOF, FORCE_CRCERR, EN_UTM_SPDUP, ATPG_ENI;
output TXVALID, DIS_STUFF, TXCRCEN, TXCRCRST, USBPOP, PKTXEND, TXCRCPHASE, 
    SOF_DISCONN, TURNCNT_EN;
    wire TXBCNT438_7, TX_HOSTDAT1397_6, TURNCNT_EN488, MACDATA388_17, 
        SOF_DISCONN_T, TX_HOSTDAT_N1352_2, MACDATA388_30, POPCNT1095_3, 
        SPAREO6, TXBCNT446_8, MACDATA_31, TXCRC5_T, HOSTTMP_5, MACDATA_16, 
        PKTXEND_4T, TX_HOSTDAT_1, MACDATA388_4, TURN_CNT543_3, POPCNT_7, 
        TXSM350_6, HOSTD978_2, MACDATA_7, POPCNT_10, MACDATA388_39, 
        SOF_DISCONN_P3, MACDATA_23, TXBCNT446_1, EOPCNT874_0, MACDATA_38, 
        TX_HOSTDAT_N1348_7, MACDATA388_22, POPCNT1087_7, POPCNT1087_10, 
        HOSTTMP1039_7, TEST_STATE310, PKTXEND_2T, POPCNT_9, POPCNT1087_0, 
        TURN_CNT535_3, HOSTTMP1039_0, PKTXEND_T, TURN_CNT_2, MACDATA_18, 
        MACDATA388_25, TX_HOSTDAT_N1348_0, SPAREO0_, MACDATA388_19, SPAREO8, 
        MACDATA_24, TXBCNT446_6, BYTECNT_1, TXSTART_T584, TXBCNT438_9, 
        MACDATA_0, n_3829, BYTECNT836_3, POPCNT1087_9, TXSM350_1, HOSTD978_5, 
        POPCNT_0, TX_HOSTDAT_6, MACDATA388_3, MACDATA_11, HOSTTMP_2, TXSM_0, 
        MACDATA_36, MACDATA388_37, TX_HOSTDAT_N1352_5, MACDATA388_10, SPAREO1, 
        MACDATA_9, POPCNT1095_4, val1280_1, TX_HOSTDAT1397_1, TXBCNT438_0, 
        TXBCNT438_8, MACDATA_1, BYTECNT836_2, MACDATA388_18, SPAREO9, 
        TXBCNT446_7, MACDATA_25, MACDATA_19, TURN_CNT_3, MACDATA388_24, 
        TX_HOSTDAT_N1348_1, POPCNT_8, POPCNT1087_1, HOSTTMP1039_1, 
        TURN_CNT535_2, START621, MACDATA_8, TXBCNT438_1, TX_HOSTDAT1397_0, 
        MACDATA388_36, TX_HOSTDAT_N1352_4, MACDATA388_11, SPAREO0, 
        POPCNT1095_5, TXRDY, HOSTTMP_3, MACDATA_10, TXSM_1, MACDATA_37, 
        BYTECNT_0, TXSM350_0, HOSTD978_4, POPCNT_1, POPCNT1087_8, TX_HOSTDAT_7, 
        MACDATA388_2, MACDATA388_5, TURN_CNT543_2, TEST_FLAG1306, POPCNT_6, 
        HOSTD978_3, TXSM_6, MACDATA_30, MACDATA_17, HOSTTMP_4, MACDATA388_16, 
        TXBCNT446_10, TX_HOSTDAT_N1352_3, MACDATA388_31, POPCNT1095_2, SPAREO7, 
        TXBCNT446_9, TX_HOSTDAT1397_7, TXBCNT438_6, USBPOP1137, POPCNT1087_6, 
        HOSTTMP1039_6, POPCNT1095_10, TEST_FLAG, TXCRC16_T, EOPCNT874_1, 
        MACDATA_39, EOPCNT_4, TX_HOSTDAT_N1348_6, MACDATA388_23, MACDATA388_38, 
        SOF_DISCONN_P2, MACDATA_22, TXBCNT446_0, MACDATA_6, TXBCNT438_4, 
        TX_HOSTDAT1397_5, n_2892, MACDATA_29, POPCNT1095_0, SPAREO5, 
        TX_HOSTDAT_N1352_1, MACDATA388_33, MACDATA388_14, MACDATA388_28, 
        MACDATA_15, HOSTTMP_6, TXSM_4, MACDATA_32, n_2889, POPCNT_4, TXSM350_5, 
        HOSTD978_1, TX_HOSTDAT_2, MACDATA388_7, TURN_CNT543_0, TXBCNTRST_, 
        MACDATA_4, POPCNT1095_9, MACDATA_20, TXBCNT446_2, SOF_CHK_COND, 
        TX_HOSTDAT_N1348_4, MACDATA388_21, EOPCNT874_3, n_4084, HOSTTMP1039_4, 
        POPCNT1087_4, TURN_CNT535_0, HOSTTMP1039_3, POPCNT1087_3, MACDATA388_9, 
        MACDATA388_26, TX_HOSTDAT_N1348_3, TURN_CNT_1, BYTECNTRST_, n_4083, 
        EOPCNT874_4, MACDATA_27, TXBCNT446_5, START, BYTECNT836_0, MACDATA_3, 
        BYTECNT_2, TX_HOSTDAT_5, MACDATA388_0, TXSM350_2, HOSTD978_6, POPCNT_3, 
        TXSM_3, MACDATA_35, HOSTTMP_1, MACDATA_12, SPAREO2, POPCNT1095_7, 
        SOF_DISCONN_P, MACDATA388_13, MACDATA388_34, TX_HOSTDAT_N1352_6, 
        TX_HOSTDAT1397_2, TXBCNT438_3, BYTECNT836_1, MACDATA_2, TXCRC5_T732, 
        TXBCNT446_4, MACDATA_26, EOPCNT_0, MACDATA388_27, TX_HOSTDAT_N1348_2, 
        TURN_CNT_0, TURN_CNT535_1, HOSTTMP1039_2, NXTISSYNC, POPCNT1087_2, 
        MACDATA388_8, PKTXEND_3T, TXBCNT438_2, TX_HOSTDAT1397_3, SPAREO3, 
        POPCNT1095_6, SPAREO1_, MACDATA388_12, MACDATA388_35, 
        TX_HOSTDAT_N1352_7, TXSM_2, MACDATA_34, MACDATA_13, BYTECNT_3, 
        TX_HOSTDAT_4, MACDATA388_1, TXSM350_3, HOSTD978_7, POPCNT_2, POPCNT_5, 
        TXSM350_4, HOSTD978_0, TX_HOSTDAT_3, MACDATA388_6, TURN_CNT543_1, 
        MACDATA388_29, val810_1, HOSTTMP_7, MACDATA_14, MACDATA_33, MACDATA_28, 
        POPCNT1095_1, SPAREO4, MACDATA388_32, MACDATA388_15, TXBCNT438_10, 
        TX_HOSTDAT1397_4, TXSTART_T, TXBCNT438_5, HOSTTMP1039_5, POPCNT1087_5, 
        TX_HOSTDAT_N1348_5, MACDATA388_20, EOPCNT874_2, POPCNT1095_8, 
        MACDATA_21, TXBCNT446_3, TXVALID658, MACDATA_5, n1685, n1917, n1918, 
        n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
        n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
        n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
        n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
        n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, 
        n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
        n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, 
        n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
        n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
        n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, 
        n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
        n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, 
        n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, 
        n2050, n2051, n2052, n2053, n2054, n2055, add_272_carry_8, 
        add_272_carry_6, add_272_carry_7, add_272_carry_9, add_272_carry_2, 
        add_272_carry_5, add_272_carry_10, add_272_carry_4, add_272_carry_3, 
        add_327_carry_2, add_327_carry_3, add_498_carry_8, add_498_carry_6, 
        add_498_carry_7, add_498_carry_9, add_498_carry_2, add_498_carry_5, 
        add_498_carry_10, add_498_carry_4, add_498_carry_3, add_549_carry_6, 
        add_549_carry_7, add_549_carry_2, add_549_carry_5, add_549_carry_4, 
        add_549_carry_3, sub_551_carry_1, sub_551_carry_7, sub_551_carry_6, 
        sub_551_carry_5, sub_551_carry_2, sub_551_carry_4, sub_551_carry_3, 
        n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, 
        n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, 
        n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, 
        n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, 
        n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, 
        n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, 
        n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, 
        n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, 
        n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, 
        n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, 
        n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, 
        n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, 
        n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, 
        n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, 
        n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, 
        n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, 
        n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, 
        n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, 
        n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, 
        n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, 
        n2256, n2257, n2258, n2259;
    zaoi211b SPARE672 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE675 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zoai21b SPARE674 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE673 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zivb SPARE678 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE671 ( .CK(CLK60M), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    znr3b SPARE676 ( .A(SPAREO2), .B(NXTISSYNC), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE677 ( .A(SPAREO4), .Y(SPAREO5) );
    znd3b SPARE679 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE670 ( .CK(CLK60M), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zxo2b U672 ( .A(n1965), .B(POPCNT_6), .Y(n2036) );
    zxo2b U673 ( .A(TXBCNT[4]), .B(n1946), .Y(n1917) );
    zxo2b U674 ( .A(n1953), .B(TXBCNT[5]), .Y(n1924) );
    zbfp U675 ( .A(MAXLEN[2]), .Y(n1951) );
    zbfp U676 ( .A(MAXLEN[3]), .Y(n1963) );
    zxo2d U677 ( .A(TXBCNT[0]), .B(n1962), .Y(n1918) );
    zxo2d U678 ( .A(n1952), .B(TXBCNT[10]), .Y(n1919) );
    zxo2d U679 ( .A(TXBCNT[8]), .B(n1956), .Y(n1920) );
    zxo2d U680 ( .A(TXBCNT[9]), .B(n1966), .Y(n1921) );
    zxo2d U681 ( .A(n1951), .B(TXBCNT[2]), .Y(n1922) );
    zxo2d U682 ( .A(TXBCNT[3]), .B(n1963), .Y(n1923) );
    zor2b U683 ( .A(TXVALID), .B(n2057), .Y(n_4083) );
    zan2b U684 ( .A(TXSM_1), .B(n2124), .Y(n2123) );
    znr2b U685 ( .A(n2124), .B(n2151), .Y(n1986) );
    znd2b U686 ( .A(n1974), .B(n2151), .Y(n2159) );
    zivb U687 ( .A(n2124), .Y(n1974) );
    znd2b U688 ( .A(n2157), .B(n2065), .Y(n2124) );
    zan3b U689 ( .A(n2151), .B(TXSM_4), .C(n2157), .Y(n2022) );
    znr2b U690 ( .A(n2137), .B(BYTECNT_1), .Y(n1984) );
    znd2b U691 ( .A(n2012), .B(n2126), .Y(n1983) );
    znr2b U692 ( .A(HANDSHK), .B(TOKEN), .Y(n2049) );
    zxo2b U693 ( .A(POPCNT_0), .B(n1962), .Y(n2014) );
    zxo2b U694 ( .A(POPCNT_7), .B(MAXLEN[7]), .Y(n2039) );
    zxo2b U695 ( .A(POPCNT_4), .B(n1946), .Y(n2038) );
    zao22b U696 ( .A(n1930), .B(CRC[4]), .C(ADRENDPS[15]), .D(n1927), .Y(n2230
        ) );
    zao22b U697 ( .A(n1930), .B(CRC[3]), .C(ADRENDPS[14]), .D(n1927), .Y(n2231
        ) );
    zao22b U698 ( .A(n1930), .B(CRC[2]), .C(ADRENDPS[13]), .D(n1927), .Y(n2232
        ) );
    zao22b U699 ( .A(n1930), .B(CRC[1]), .C(ADRENDPS[12]), .D(n1927), .Y(n2233
        ) );
    zao22b U700 ( .A(n1930), .B(CRC[0]), .C(ADRENDPS[11]), .D(n1927), .Y(n2234
        ) );
    zivb U701 ( .A(SPLIT), .Y(n1980) );
    zan2b U702 ( .A(MACDATA_10), .B(n2241), .Y(n2148) );
    zan2b U703 ( .A(MACDATA_8), .B(n1942), .Y(n2141) );
    zan2b U704 ( .A(ADRENDPS[7]), .B(n1934), .Y(n2142) );
    znd2b U705 ( .A(n1993), .B(n1994), .Y(n2206) );
    zmux21lb U706 ( .A(n1940), .B(n1941), .S(CRC[7]), .Y(n1993) );
    zan2b U707 ( .A(ADRENDPS[6]), .B(n1934), .Y(n2143) );
    znd2b U708 ( .A(n1995), .B(n1996), .Y(n2209) );
    zmux21lb U709 ( .A(n1940), .B(n1941), .S(CRC[6]), .Y(n1995) );
    zan2b U710 ( .A(ADRENDPS[5]), .B(n1934), .Y(n2144) );
    znd2b U711 ( .A(n1997), .B(n1998), .Y(n2212) );
    zmux21lb U712 ( .A(n1940), .B(n1941), .S(CRC[5]), .Y(n1997) );
    zan2b U713 ( .A(ADRENDPS[4]), .B(n1934), .Y(n2145) );
    znd2b U714 ( .A(n1999), .B(n2000), .Y(n2215) );
    zmux21lb U715 ( .A(n1940), .B(n1941), .S(CRC[4]), .Y(n1999) );
    zan2b U716 ( .A(ADRENDPS[3]), .B(n1934), .Y(n2146) );
    znd2b U717 ( .A(n2001), .B(n2002), .Y(n2218) );
    zmux21lb U718 ( .A(n1940), .B(n1941), .S(CRC[3]), .Y(n2001) );
    zan2b U719 ( .A(ADRENDPS[2]), .B(n1934), .Y(n2147) );
    znd2b U720 ( .A(n2003), .B(n2004), .Y(n2221) );
    zmux21lb U721 ( .A(n1940), .B(n1941), .S(CRC[2]), .Y(n2003) );
    zan2b U722 ( .A(ADRENDPS[1]), .B(n1934), .Y(n2149) );
    znd2b U723 ( .A(n2005), .B(n2006), .Y(n2224) );
    zmux21lb U724 ( .A(n1940), .B(n1941), .S(CRC[1]), .Y(n2005) );
    zor2b U725 ( .A(n2176), .B(n2177), .Y(n2203) );
    zor2b U726 ( .A(n2236), .B(n2176), .Y(n2202) );
    zivb U727 ( .A(n2177), .Y(n2236) );
    znd2b U728 ( .A(n1970), .B(n1971), .Y(n2177) );
    zivb U729 ( .A(SL_FORCE_CRC), .Y(n1970) );
    zivb U730 ( .A(FORCE_CRCERR), .Y(n1971) );
    zcxi4b U731 ( .A(n2054), .B(n2186), .C(n1991), .D(n1992), .Y(n2226) );
    znr2b U732 ( .A(n1990), .B(n2011), .Y(n1991) );
    zivb U733 ( .A(ADRENDPS[0]), .Y(n2011) );
    zor2b U734 ( .A(TXSM_6), .B(n2167), .Y(n2171) );
    zivb U735 ( .A(n2171), .Y(n2173) );
    zivb U736 ( .A(n2178), .Y(n2174) );
    zor2b sub_551_U1_B_6 ( .A(TX_HOSTDAT_6), .B(sub_551_carry_6), .Y(
        sub_551_carry_7) );
    zor2b sub_551_U1_B_5 ( .A(TX_HOSTDAT_5), .B(sub_551_carry_5), .Y(
        sub_551_carry_6) );
    zor2b sub_551_U1_B_4 ( .A(TX_HOSTDAT_4), .B(sub_551_carry_4), .Y(
        sub_551_carry_5) );
    zor2b sub_551_U1_B_3 ( .A(TX_HOSTDAT_3), .B(sub_551_carry_3), .Y(
        sub_551_carry_4) );
    zor2b sub_551_U1_B_2 ( .A(TX_HOSTDAT_2), .B(sub_551_carry_2), .Y(
        sub_551_carry_3) );
    zor2b sub_551_U1_B_1 ( .A(TX_HOSTDAT_1), .B(sub_551_carry_1), .Y(
        sub_551_carry_2) );
    zaoi2x4b U737 ( .A(n2130), .B(n2131), .C(n1926), .D(n2132), .E(HANDSHK), 
        .F(n2133), .G(BYTECNT_1), .H(n2134), .Y(n2129) );
    zmux21lb U738 ( .A(n2077), .B(n2078), .S(SPLIT), .Y(n2130) );
    zivb U739 ( .A(n2137), .Y(n2134) );
    znd3b U740 ( .A(TXCRCPHASE), .B(n1972), .C(n2155), .Y(n2137) );
    zxo2b U741 ( .A(TURN_CNT_0), .B(TURN_PARM[0]), .Y(n2197) );
    zxo2b U742 ( .A(TURN_CNT_2), .B(TURN_PARM[2]), .Y(n2196) );
    zxo2b U743 ( .A(TURN_CNT_3), .B(TURN_PARM[3]), .Y(n2199) );
    zxo2b U744 ( .A(TURN_CNT_1), .B(TURN_PARM[1]), .Y(n2198) );
    zoa22b U745 ( .A(BYTECNT_3), .B(n2127), .C(n2136), .D(n2057), .Y(n2135) );
    znd2b U746 ( .A(n2056), .B(BYTECNT_3), .Y(n2050) );
    znd2b U747 ( .A(n1968), .B(TXVALID), .Y(n2021) );
    zan3b U748 ( .A(n1926), .B(n2122), .C(n1968), .Y(n2121) );
    zor2b U749 ( .A(EOPCNT_4), .B(n2128), .Y(n2122) );
    zivb U750 ( .A(n2122), .Y(n2132) );
    zivb U751 ( .A(n2136), .Y(n2229) );
    zxo2b U752 ( .A(n2154), .B(n2155), .Y(n2153) );
    znd2b U753 ( .A(n2067), .B(n1972), .Y(n2154) );
    zivb U754 ( .A(n2127), .Y(n2048) );
    znd2b U755 ( .A(n1986), .B(n1987), .Y(n2127) );
    zmux21lb U756 ( .A(BYTECNT_2), .B(BYTECNT_3), .S(SPLIT), .Y(n2053) );
    zor2b U757 ( .A(TXVALID), .B(START), .Y(n1977) );
    znr2b U758 ( .A(n2154), .B(n2125), .Y(n1975) );
    zivb U759 ( .A(n2160), .Y(n1976) );
    znd2b U760 ( .A(n2158), .B(n1985), .Y(n2160) );
    zivb U761 ( .A(n2159), .Y(n1985) );
    znd2b U762 ( .A(n1987), .B(n2022), .Y(n2012) );
    zivb U763 ( .A(n2156), .Y(n1987) );
    zor2b U764 ( .A(TXSM_1), .B(n2152), .Y(n2235) );
    znd2b U765 ( .A(DIS_STUFF), .B(n1969), .Y(n2120) );
    zao2x4b U766 ( .A(sub_551_carry_1), .B(n2069), .C(SL_TXFIXDATA[0]), .D(
        n2070), .E(TX_HOSTDAT_N1348_0), .F(n2071), .G(TX_HOSTDAT_N1348_0), .H(
        n2072), .Y(TX_HOSTDAT1397_0) );
    zor2b U767 ( .A(MACDATA_39), .B(n2115), .Y(MACDATA388_39) );
    zor2b U768 ( .A(MACDATA_38), .B(n2115), .Y(MACDATA388_38) );
    zor2b U769 ( .A(MACDATA_37), .B(n2115), .Y(MACDATA388_37) );
    zor2b U770 ( .A(MACDATA_36), .B(n2115), .Y(MACDATA388_36) );
    zor2b U771 ( .A(MACDATA_35), .B(n2115), .Y(MACDATA388_35) );
    zor2b U772 ( .A(MACDATA_34), .B(n2115), .Y(MACDATA388_34) );
    zor2b U773 ( .A(MACDATA_33), .B(n2115), .Y(MACDATA388_33) );
    zor2b U774 ( .A(MACDATA_32), .B(n2115), .Y(MACDATA388_32) );
    zao21b U775 ( .A(MACDATA_39), .B(n2240), .C(n2114), .Y(MACDATA388_31) );
    zan2b U776 ( .A(MACDATA_29), .B(n1942), .Y(n2112) );
    zan2b U777 ( .A(MACDATA_27), .B(n1942), .Y(n2110) );
    zan2b U778 ( .A(MACDATA_25), .B(n2241), .Y(n2108) );
    zao22b U779 ( .A(n1927), .B(CRC[4]), .C(MACDATA_23), .D(n2241), .Y(n2106)
         );
    zao22b U780 ( .A(CRC[2]), .B(n1927), .C(MACDATA_21), .D(n2241), .Y(n2104)
         );
    zao22b U781 ( .A(CRC[0]), .B(n1927), .C(MACDATA_19), .D(n1942), .Y(n2102)
         );
    zao22b U782 ( .A(ADRENDPS[16]), .B(n1927), .C(MACDATA_16), .D(n1942), .Y(
        n2098) );
    zmux21lb U783 ( .A(n2202), .B(n2203), .S(CRC[15]), .Y(n2096) );
    zmux21lb U784 ( .A(n2202), .B(n2203), .S(CRC[14]), .Y(n2094) );
    zmux21lb U785 ( .A(n2202), .B(n2203), .S(CRC[13]), .Y(n2092) );
    zmux21lb U786 ( .A(n2202), .B(n2203), .S(CRC[12]), .Y(n2090) );
    zmux21lb U787 ( .A(n2202), .B(n2203), .S(CRC[11]), .Y(n2088) );
    zmux21lb U788 ( .A(n2202), .B(n2203), .S(CRC[10]), .Y(n2087) );
    zivb U789 ( .A(n2237), .Y(n2242) );
    zmux21lb U790 ( .A(n2202), .B(n2203), .S(CRC[9]), .Y(n2085) );
    zivb U791 ( .A(n2237), .Y(n2099) );
    zmux21lb U792 ( .A(n2202), .B(n2203), .S(CRC[8]), .Y(n2083) );
    zmux21hb U793 ( .A(n2204), .B(MACDATA_7), .S(n1942), .Y(MACDATA388_7) );
    zmux21hb U794 ( .A(n2211), .B(MACDATA_5), .S(n2241), .Y(MACDATA388_5) );
    zmux21hb U795 ( .A(n2217), .B(MACDATA_3), .S(n1942), .Y(MACDATA388_3) );
    zmux21hb U796 ( .A(n2223), .B(MACDATA_1), .S(n2241), .Y(MACDATA388_1) );
    zivb U797 ( .A(n2172), .Y(n2205) );
    zivb U798 ( .A(n2115), .Y(n2241) );
    zivb U799 ( .A(n2021), .Y(n2056) );
    zivb U800 ( .A(n2235), .Y(NXTISSYNC) );
    zcx3b U801 ( .A(MACDATA_8), .B(n2079), .C(n2080), .D(n2081), .Y(
        MACDATA388_0) );
    zivb U802 ( .A(n2175), .Y(n2079) );
    zmux21lb U803 ( .A(n2239), .B(n2238), .S(CRC[0]), .Y(n2081) );
    zivb U804 ( .A(n2202), .Y(n2239) );
    zivb U805 ( .A(n2203), .Y(n2238) );
    zivb U806 ( .A(n2175), .Y(n2240) );
    zxo2b U807 ( .A(add_272_carry_10), .B(TXBCNT[10]), .Y(TXBCNT438_10) );
    zhadrb add_272_U1_1_9 ( .A(TXBCNT[9]), .B(add_272_carry_9), .CO(
        add_272_carry_10), .S(TXBCNT438_9) );
    zhadrb add_272_U1_1_8 ( .A(TXBCNT[8]), .B(add_272_carry_8), .CO(
        add_272_carry_9), .S(TXBCNT438_8) );
    zhadrb add_272_U1_1_7 ( .A(TXBCNT[7]), .B(add_272_carry_7), .CO(
        add_272_carry_8), .S(TXBCNT438_7) );
    zhadrb add_272_U1_1_6 ( .A(TXBCNT[6]), .B(add_272_carry_6), .CO(
        add_272_carry_7), .S(TXBCNT438_6) );
    zhadrb add_272_U1_1_4 ( .A(TXBCNT[4]), .B(add_272_carry_4), .CO(
        add_272_carry_5), .S(TXBCNT438_4) );
    zhadrb add_272_U1_1_2 ( .A(TXBCNT[2]), .B(add_272_carry_2), .CO(
        add_272_carry_3), .S(TXBCNT438_2) );
    zhadrb add_272_U1_1_1 ( .A(TXBCNT[1]), .B(TXBCNT[0]), .CO(add_272_carry_2), 
        .S(TXBCNT438_1) );
    zan2b U808 ( .A(TURNCNT_EN), .B(TURN_CNT535_3), .Y(TURN_CNT543_3) );
    zxo2b U809 ( .A(add_327_carry_3), .B(TURN_CNT_3), .Y(TURN_CNT535_3) );
    zan2b U810 ( .A(TURN_CNT535_2), .B(TURNCNT_EN), .Y(TURN_CNT543_2) );
    zhadrb add_327_U1_1_2 ( .A(TURN_CNT_2), .B(add_327_carry_2), .CO(
        add_327_carry_3), .S(TURN_CNT535_2) );
    zan2b U811 ( .A(TURN_CNT535_1), .B(TURNCNT_EN), .Y(TURN_CNT543_1) );
    zhadrb add_327_U1_1_1 ( .A(TURN_CNT_1), .B(TURN_CNT_0), .CO(
        add_327_carry_2), .S(TURN_CNT535_1) );
    zan2b U812 ( .A(TURN_CNT535_0), .B(TURNCNT_EN), .Y(TURN_CNT543_0) );
    zivb U813 ( .A(SL_TXDATASEL[2]), .Y(n2195) );
    zmux21lb U814 ( .A(n2179), .B(n2187), .S(TXRDY), .Y(HOSTTMP1039_7) );
    zmux21lb U815 ( .A(n2180), .B(n2188), .S(TXRDY), .Y(HOSTTMP1039_6) );
    zmux21lb U816 ( .A(n2181), .B(n2189), .S(TXRDY), .Y(HOSTTMP1039_5) );
    zmux21lb U817 ( .A(n2182), .B(n2190), .S(TXRDY), .Y(HOSTTMP1039_4) );
    zmux21lb U818 ( .A(n2183), .B(n2191), .S(TXRDY), .Y(HOSTTMP1039_3) );
    zmux21lb U819 ( .A(n2184), .B(n2192), .S(TXRDY), .Y(HOSTTMP1039_2) );
    zmux21lb U820 ( .A(n2185), .B(n2193), .S(TXRDY), .Y(HOSTTMP1039_1) );
    zmux21lb U821 ( .A(n2186), .B(n2194), .S(TXRDY), .Y(HOSTTMP1039_0) );
    zxo2b U822 ( .A(add_498_carry_10), .B(POPCNT_10), .Y(POPCNT1087_10) );
    zhadrb add_498_U1_1_9 ( .A(POPCNT_9), .B(add_498_carry_9), .CO(
        add_498_carry_10), .S(POPCNT1087_9) );
    zhadrb add_498_U1_1_8 ( .A(POPCNT_8), .B(add_498_carry_8), .CO(
        add_498_carry_9), .S(POPCNT1087_8) );
    zhadrb add_498_U1_1_7 ( .A(POPCNT_7), .B(add_498_carry_7), .CO(
        add_498_carry_8), .S(POPCNT1087_7) );
    zhadrb add_498_U1_1_6 ( .A(POPCNT_6), .B(add_498_carry_6), .CO(
        add_498_carry_7), .S(POPCNT1087_6) );
    zhadrb add_498_U1_1_5 ( .A(POPCNT_5), .B(add_498_carry_5), .CO(
        add_498_carry_6), .S(POPCNT1087_5) );
    zhadrb add_498_U1_1_4 ( .A(POPCNT_4), .B(add_498_carry_4), .CO(
        add_498_carry_5), .S(POPCNT1087_4) );
    zhadrb add_498_U1_1_3 ( .A(POPCNT_3), .B(add_498_carry_3), .CO(
        add_498_carry_4), .S(POPCNT1087_3) );
    zhadrb add_498_U1_1_2 ( .A(POPCNT_2), .B(add_498_carry_2), .CO(
        add_498_carry_3), .S(POPCNT1087_2) );
    zhadrb add_498_U1_1_1 ( .A(POPCNT_1), .B(POPCNT_0), .CO(add_498_carry_2), 
        .S(POPCNT1087_1) );
    zao2x4b U823 ( .A(n2069), .B(TX_HOSTDAT_7), .C(SL_TXFIXDATA[7]), .D(n2070), 
        .E(TX_HOSTDAT_N1348_7), .F(n2071), .G(TX_HOSTDAT_N1352_7), .H(n2072), 
        .Y(TX_HOSTDAT1397_7) );
    zxo2b U824 ( .A(add_549_carry_7), .B(TX_HOSTDAT_7), .Y(TX_HOSTDAT_N1348_7)
         );
    zxn2b sub_551_U1_A_7 ( .A(TX_HOSTDAT_7), .B(sub_551_carry_7), .Y(
        TX_HOSTDAT_N1352_7) );
    zao2x4b U825 ( .A(TX_HOSTDAT_6), .B(n2069), .C(SL_TXFIXDATA[6]), .D(n2070), 
        .E(TX_HOSTDAT_N1348_6), .F(n2071), .G(TX_HOSTDAT_N1352_6), .H(n2072), 
        .Y(TX_HOSTDAT1397_6) );
    zhadrb add_549_U1_1_6 ( .A(TX_HOSTDAT_6), .B(add_549_carry_6), .CO(
        add_549_carry_7), .S(TX_HOSTDAT_N1348_6) );
    zxn2b sub_551_U1_A_6 ( .A(TX_HOSTDAT_6), .B(sub_551_carry_6), .Y(
        TX_HOSTDAT_N1352_6) );
    zao2x4b U826 ( .A(TX_HOSTDAT_5), .B(n2069), .C(SL_TXFIXDATA[5]), .D(n2070), 
        .E(TX_HOSTDAT_N1348_5), .F(n2071), .G(TX_HOSTDAT_N1352_5), .H(n2072), 
        .Y(TX_HOSTDAT1397_5) );
    zhadrb add_549_U1_1_5 ( .A(TX_HOSTDAT_5), .B(add_549_carry_5), .CO(
        add_549_carry_6), .S(TX_HOSTDAT_N1348_5) );
    zxn2b sub_551_U1_A_5 ( .A(TX_HOSTDAT_5), .B(sub_551_carry_5), .Y(
        TX_HOSTDAT_N1352_5) );
    zao2x4b U827 ( .A(TX_HOSTDAT_4), .B(n2069), .C(SL_TXFIXDATA[4]), .D(n2070), 
        .E(TX_HOSTDAT_N1348_4), .F(n2071), .G(TX_HOSTDAT_N1352_4), .H(n2072), 
        .Y(TX_HOSTDAT1397_4) );
    zhadrb add_549_U1_1_4 ( .A(TX_HOSTDAT_4), .B(add_549_carry_4), .CO(
        add_549_carry_5), .S(TX_HOSTDAT_N1348_4) );
    zxn2b sub_551_U1_A_4 ( .A(TX_HOSTDAT_4), .B(sub_551_carry_4), .Y(
        TX_HOSTDAT_N1352_4) );
    zao2x4b U828 ( .A(TX_HOSTDAT_3), .B(n2069), .C(SL_TXFIXDATA[3]), .D(n2070), 
        .E(TX_HOSTDAT_N1348_3), .F(n2071), .G(TX_HOSTDAT_N1352_3), .H(n2072), 
        .Y(TX_HOSTDAT1397_3) );
    zhadrb add_549_U1_1_3 ( .A(TX_HOSTDAT_3), .B(add_549_carry_3), .CO(
        add_549_carry_4), .S(TX_HOSTDAT_N1348_3) );
    zxn2b sub_551_U1_A_3 ( .A(TX_HOSTDAT_3), .B(sub_551_carry_3), .Y(
        TX_HOSTDAT_N1352_3) );
    zao2x4b U829 ( .A(TX_HOSTDAT_2), .B(n2069), .C(SL_TXFIXDATA[2]), .D(n2070), 
        .E(TX_HOSTDAT_N1348_2), .F(n2071), .G(TX_HOSTDAT_N1352_2), .H(n2072), 
        .Y(TX_HOSTDAT1397_2) );
    zhadrb add_549_U1_1_2 ( .A(TX_HOSTDAT_2), .B(add_549_carry_2), .CO(
        add_549_carry_3), .S(TX_HOSTDAT_N1348_2) );
    zxn2b sub_551_U1_A_2 ( .A(TX_HOSTDAT_2), .B(sub_551_carry_2), .Y(
        TX_HOSTDAT_N1352_2) );
    zivd U830 ( .A(n2163), .Y(n2072) );
    zao2x4b U831 ( .A(TX_HOSTDAT_1), .B(n2069), .C(SL_TXFIXDATA[1]), .D(n2070), 
        .E(TX_HOSTDAT_N1348_1), .F(n2071), .G(TX_HOSTDAT_N1352_1), .H(n2072), 
        .Y(TX_HOSTDAT1397_1) );
    zivc U832 ( .A(n2165), .Y(n2069) );
    zhadrb add_549_U1_1_1 ( .A(TX_HOSTDAT_1), .B(sub_551_carry_1), .CO(
        add_549_carry_2), .S(TX_HOSTDAT_N1348_1) );
    zivc U833 ( .A(n2164), .Y(n2071) );
    zxn2b sub_551_U1_A_1 ( .A(TX_HOSTDAT_1), .B(sub_551_carry_1), .Y(
        TX_HOSTDAT_N1352_1) );
    zivb U834 ( .A(SL_TXDATASEL[0]), .Y(n2162) );
    zor2b U835 ( .A(n2166), .B(n2129), .Y(n2167) );
    zor2b U836 ( .A(n2166), .B(n2135), .Y(n2152) );
    zivb U837 ( .A(n1977), .Y(n2166) );
    zmux21hb U838 ( .A(TXCRC16_T), .B(TXCRC5_T), .S(TOKEN), .Y(val810_1) );
    zan2b U839 ( .A(n1933), .B(TXSTART_T), .Y(START621) );
    zmux21hb U840 ( .A(PKTXEND_3T), .B(n1925), .S(EN_UTM_SPDUP), .Y(val1280_1)
         );
    znr5b U841 ( .A(n2058), .B(TEST_J), .C(TEST_PACKET), .D(TEST_EYE), .E(
        TEST_K), .Y(SOF_CHK_COND) );
    zivb U842 ( .A(TXSOF), .Y(n2128) );
    zivb U843 ( .A(n2120), .Y(n2150) );
    zivb U844 ( .A(n1981), .Y(n2117) );
    zoai21b U845 ( .A(n1933), .B(n2059), .C(n2060), .Y(TXSTART_T584) );
    zivd U846 ( .A(TXSTART), .Y(n2060) );
    zan3b U847 ( .A(n1968), .B(TXSM_1), .C(n2061), .Y(TXCRC5_T732) );
    zivb U848 ( .A(n2064), .Y(n1979) );
    zan2b U849 ( .A(SOF_DISCONN_P2), .B(SOF_DISCONN_P3), .Y(n2062) );
    zivb U850 ( .A(DIS_STUFF), .Y(n2118) );
    zmux21hb U851 ( .A(MACDATA_0), .B(n_2892), .S(n1685), .Y(DATA_TX[0]) );
    zmux21hb U852 ( .A(MACDATA_1), .B(n_2889), .S(n1685), .Y(DATA_TX[1]) );
    zmux21hb U853 ( .A(MACDATA_2), .B(n_2889), .S(n1685), .Y(DATA_TX[2]) );
    zmux21hb U854 ( .A(MACDATA_3), .B(n_2889), .S(n1685), .Y(DATA_TX[3]) );
    zmux21hb U855 ( .A(MACDATA_4), .B(n_2889), .S(n1685), .Y(DATA_TX[4]) );
    zmux21hb U856 ( .A(MACDATA_5), .B(n_2889), .S(n1685), .Y(DATA_TX[5]) );
    zmux21hb U857 ( .A(MACDATA_6), .B(n_2889), .S(n1685), .Y(DATA_TX[6]) );
    zmux21hb U858 ( .A(MACDATA_7), .B(n_2889), .S(n1685), .Y(DATA_TX[7]) );
    zivb U859 ( .A(TEST_EYE), .Y(n_2889) );
    zivb U860 ( .A(BYTECNT_3), .Y(n2078) );
    zdffqrb MACDATA_reg_39 ( .CK(CLK60M), .D(MACDATA388_39), .R(TRST_), .Q(
        MACDATA_39) );
    zdffqrb MACDATA_reg_38 ( .CK(CLK60M), .D(MACDATA388_38), .R(TRST_), .Q(
        MACDATA_38) );
    zdffqrb MACDATA_reg_37 ( .CK(CLK60M), .D(MACDATA388_37), .R(TRST_), .Q(
        MACDATA_37) );
    zdffqrb MACDATA_reg_36 ( .CK(CLK60M), .D(MACDATA388_36), .R(TRST_), .Q(
        MACDATA_36) );
    zdffqrb MACDATA_reg_35 ( .CK(CLK60M), .D(MACDATA388_35), .R(TRST_), .Q(
        MACDATA_35) );
    zdffqrb MACDATA_reg_34 ( .CK(CLK60M), .D(MACDATA388_34), .R(TRST_), .Q(
        MACDATA_34) );
    zdffqrb MACDATA_reg_33 ( .CK(CLK60M), .D(MACDATA388_33), .R(TRST_), .Q(
        MACDATA_33) );
    zdffqrb MACDATA_reg_32 ( .CK(CLK60M), .D(MACDATA388_32), .R(TRST_), .Q(
        MACDATA_32) );
    zdffqrb MACDATA_reg_31 ( .CK(CLK60M), .D(MACDATA388_31), .R(TRST_), .Q(
        MACDATA_31) );
    zdffqrb MACDATA_reg_30 ( .CK(CLK60M), .D(MACDATA388_30), .R(TRST_), .Q(
        MACDATA_30) );
    zdffqrb MACDATA_reg_29 ( .CK(CLK60M), .D(MACDATA388_29), .R(TRST_), .Q(
        MACDATA_29) );
    zdffqrb MACDATA_reg_28 ( .CK(CLK60M), .D(MACDATA388_28), .R(TRST_), .Q(
        MACDATA_28) );
    zdffqrb MACDATA_reg_27 ( .CK(CLK60M), .D(MACDATA388_27), .R(TRST_), .Q(
        MACDATA_27) );
    zdffqrb MACDATA_reg_26 ( .CK(CLK60M), .D(MACDATA388_26), .R(TRST_), .Q(
        MACDATA_26) );
    zdffqrb MACDATA_reg_25 ( .CK(CLK60M), .D(MACDATA388_25), .R(TRST_), .Q(
        MACDATA_25) );
    zdffqrb MACDATA_reg_24 ( .CK(CLK60M), .D(MACDATA388_24), .R(TRST_), .Q(
        MACDATA_24) );
    zdffqrb MACDATA_reg_23 ( .CK(CLK60M), .D(MACDATA388_23), .R(TRST_), .Q(
        MACDATA_23) );
    zdffqrb MACDATA_reg_22 ( .CK(CLK60M), .D(MACDATA388_22), .R(TRST_), .Q(
        MACDATA_22) );
    zdffqrb MACDATA_reg_21 ( .CK(CLK60M), .D(MACDATA388_21), .R(TRST_), .Q(
        MACDATA_21) );
    zdffqrb MACDATA_reg_20 ( .CK(CLK60M), .D(MACDATA388_20), .R(TRST_), .Q(
        MACDATA_20) );
    zdffqrb MACDATA_reg_19 ( .CK(CLK60M), .D(MACDATA388_19), .R(TRST_), .Q(
        MACDATA_19) );
    zdffqrb MACDATA_reg_18 ( .CK(CLK60M), .D(MACDATA388_18), .R(TRST_), .Q(
        MACDATA_18) );
    zdffqrb MACDATA_reg_17 ( .CK(CLK60M), .D(MACDATA388_17), .R(TRST_), .Q(
        MACDATA_17) );
    zdffqrb MACDATA_reg_16 ( .CK(CLK60M), .D(MACDATA388_16), .R(TRST_), .Q(
        MACDATA_16) );
    zdffqrb MACDATA_reg_15 ( .CK(CLK60M), .D(MACDATA388_15), .R(TRST_), .Q(
        MACDATA_15) );
    zdffqrb MACDATA_reg_14 ( .CK(CLK60M), .D(MACDATA388_14), .R(TRST_), .Q(
        MACDATA_14) );
    zdffqrb MACDATA_reg_13 ( .CK(CLK60M), .D(MACDATA388_13), .R(TRST_), .Q(
        MACDATA_13) );
    zdffqrb MACDATA_reg_12 ( .CK(CLK60M), .D(MACDATA388_12), .R(TRST_), .Q(
        MACDATA_12) );
    zdffqrb MACDATA_reg_11 ( .CK(CLK60M), .D(MACDATA388_11), .R(TRST_), .Q(
        MACDATA_11) );
    zdffqrb MACDATA_reg_10 ( .CK(CLK60M), .D(MACDATA388_10), .R(TRST_), .Q(
        MACDATA_10) );
    zdffqrb MACDATA_reg_9 ( .CK(CLK60M), .D(MACDATA388_9), .R(TRST_), .Q(
        MACDATA_9) );
    zdffqrb MACDATA_reg_8 ( .CK(CLK60M), .D(MACDATA388_8), .R(TRST_), .Q(
        MACDATA_8) );
    zdffqrb MACDATA_reg_7 ( .CK(CLK60M), .D(MACDATA388_7), .R(TRST_), .Q(
        MACDATA_7) );
    zdffqrb MACDATA_reg_6 ( .CK(CLK60M), .D(MACDATA388_6), .R(TRST_), .Q(
        MACDATA_6) );
    zdffqrb MACDATA_reg_5 ( .CK(CLK60M), .D(MACDATA388_5), .R(TRST_), .Q(
        MACDATA_5) );
    zdffqrb MACDATA_reg_4 ( .CK(CLK60M), .D(MACDATA388_4), .R(TRST_), .Q(
        MACDATA_4) );
    zdffqrb MACDATA_reg_3 ( .CK(CLK60M), .D(MACDATA388_3), .R(TRST_), .Q(
        MACDATA_3) );
    zdffqrb MACDATA_reg_2 ( .CK(CLK60M), .D(MACDATA388_2), .R(TRST_), .Q(
        MACDATA_2) );
    zdffqrb MACDATA_reg_1 ( .CK(CLK60M), .D(MACDATA388_1), .R(TRST_), .Q(
        MACDATA_1) );
    zdffqrb MACDATA_reg_0 ( .CK(CLK60M), .D(MACDATA388_0), .R(TRST_), .Q(
        MACDATA_0) );
    zdffqrb TXBCNT_reg_10 ( .CK(CLK60M), .D(TXBCNT446_10), .R(TXBCNTRST_), .Q(
        TXBCNT[10]) );
    zdffqrb TXBCNT_reg_9 ( .CK(CLK60M), .D(TXBCNT446_9), .R(TXBCNTRST_), .Q(
        TXBCNT[9]) );
    zdffqrb TXBCNT_reg_8 ( .CK(CLK60M), .D(TXBCNT446_8), .R(TXBCNTRST_), .Q(
        TXBCNT[8]) );
    zdffqrb TXBCNT_reg_7 ( .CK(CLK60M), .D(TXBCNT446_7), .R(TXBCNTRST_), .Q(
        TXBCNT[7]) );
    zdffqrb TXBCNT_reg_6 ( .CK(CLK60M), .D(TXBCNT446_6), .R(TXBCNTRST_), .Q(
        TXBCNT[6]) );
    zdffqrb TXBCNT_reg_4 ( .CK(CLK60M), .D(TXBCNT446_4), .R(TXBCNTRST_), .Q(
        TXBCNT[4]) );
    zdffqrb TXBCNT_reg_2 ( .CK(CLK60M), .D(TXBCNT446_2), .R(TXBCNTRST_), .Q(
        TXBCNT[2]) );
    zdffqrb TXBCNT_reg_1 ( .CK(CLK60M), .D(TXBCNT446_1), .R(TXBCNTRST_), .Q(
        TXBCNT[1]) );
    zdffqrb TXBCNT_reg_0 ( .CK(CLK60M), .D(TXBCNT446_0), .R(TXBCNTRST_), .Q(
        TXBCNT[0]) );
    zivb U861 ( .A(TXBCNT[0]), .Y(TXBCNT438_0) );
    zdffqrb TURN_CNT_reg_3 ( .CK(CLK60M), .D(TURN_CNT543_3), .R(TRST_), .Q(
        TURN_CNT_3) );
    zdffqrb TURN_CNT_reg_2 ( .CK(CLK60M), .D(TURN_CNT543_2), .R(TRST_), .Q(
        TURN_CNT_2) );
    zdffqrb TURN_CNT_reg_1 ( .CK(CLK60M), .D(TURN_CNT543_1), .R(TRST_), .Q(
        TURN_CNT_1) );
    zdffqrb TURN_CNT_reg_0 ( .CK(CLK60M), .D(TURN_CNT543_0), .R(TRST_), .Q(
        TURN_CNT_0) );
    zivb U862 ( .A(TURN_CNT_0), .Y(TURN_CNT535_0) );
    zdffqrb HOSTD_reg_7 ( .CK(CLK60M), .D(HOSTD978_7), .R(STSRST_), .Q(
        TXCRCDAT[7]) );
    zivb U863 ( .A(TXCRCDAT[7]), .Y(n2187) );
    zdffqrb HOSTD_reg_6 ( .CK(CLK60M), .D(HOSTD978_6), .R(STSRST_), .Q(
        TXCRCDAT[6]) );
    zivb U864 ( .A(TXCRCDAT[6]), .Y(n2188) );
    zdffqrb HOSTD_reg_5 ( .CK(CLK60M), .D(HOSTD978_5), .R(STSRST_), .Q(
        TXCRCDAT[5]) );
    zivb U865 ( .A(TXCRCDAT[5]), .Y(n2189) );
    zdffqrb HOSTD_reg_4 ( .CK(CLK60M), .D(HOSTD978_4), .R(STSRST_), .Q(
        TXCRCDAT[4]) );
    zivb U866 ( .A(TXCRCDAT[4]), .Y(n2190) );
    zdffqrb HOSTD_reg_3 ( .CK(CLK60M), .D(HOSTD978_3), .R(STSRST_), .Q(
        TXCRCDAT[3]) );
    zivb U867 ( .A(TXCRCDAT[3]), .Y(n2191) );
    zdffqrb HOSTD_reg_2 ( .CK(CLK60M), .D(HOSTD978_2), .R(STSRST_), .Q(
        TXCRCDAT[2]) );
    zivb U868 ( .A(TXCRCDAT[2]), .Y(n2192) );
    zdffqrb HOSTD_reg_1 ( .CK(CLK60M), .D(HOSTD978_1), .R(STSRST_), .Q(
        TXCRCDAT[1]) );
    zivb U869 ( .A(TXCRCDAT[1]), .Y(n2193) );
    zdffqrb HOSTD_reg_0 ( .CK(CLK60M), .D(HOSTD978_0), .R(STSRST_), .Q(
        TXCRCDAT[0]) );
    zivb U870 ( .A(TXCRCDAT[0]), .Y(n2194) );
    zdffrb_ HOSTTMP_reg_7 ( .CK(CLK60M), .D(n2259), .R(STSRST_), .Q(HOSTTMP_7), 
        .QN(n2179) );
    zdffrb_ HOSTTMP_reg_6 ( .CK(CLK60M), .D(n2258), .R(STSRST_), .Q(HOSTTMP_6), 
        .QN(n2180) );
    zdffrb_ HOSTTMP_reg_5 ( .CK(CLK60M), .D(n2257), .R(STSRST_), .Q(HOSTTMP_5), 
        .QN(n2181) );
    zdffrb_ HOSTTMP_reg_4 ( .CK(CLK60M), .D(n2256), .R(STSRST_), .Q(HOSTTMP_4), 
        .QN(n2182) );
    zdffrb_ HOSTTMP_reg_3 ( .CK(CLK60M), .D(n2255), .R(STSRST_), .Q(HOSTTMP_3), 
        .QN(n2183) );
    zdffrb_ HOSTTMP_reg_2 ( .CK(CLK60M), .D(n2254), .R(STSRST_), .Q(HOSTTMP_2), 
        .QN(n2184) );
    zdffrb_ HOSTTMP_reg_1 ( .CK(CLK60M), .D(n2253), .R(STSRST_), .Q(HOSTTMP_1), 
        .QN(n2185) );
    zdffrb_ HOSTTMP_reg_0 ( .CK(CLK60M), .D(HOSTTMP1039_0), .R(STSRST_), .QN(
        n2186) );
    zdffqrb POPCNT_reg_10 ( .CK(CLK60M), .D(POPCNT1095_10), .R(STSRST_), .Q(
        POPCNT_10) );
    zdffqrb POPCNT_reg_9 ( .CK(CLK60M), .D(POPCNT1095_9), .R(STSRST_), .Q(
        POPCNT_9) );
    zdffqrb POPCNT_reg_8 ( .CK(CLK60M), .D(POPCNT1095_8), .R(STSRST_), .Q(
        POPCNT_8) );
    zdffqrb POPCNT_reg_7 ( .CK(CLK60M), .D(POPCNT1095_7), .R(STSRST_), .Q(
        POPCNT_7) );
    zdffqrb POPCNT_reg_6 ( .CK(CLK60M), .D(POPCNT1095_6), .R(STSRST_), .Q(
        POPCNT_6) );
    zdffqrb POPCNT_reg_5 ( .CK(CLK60M), .D(POPCNT1095_5), .R(STSRST_), .Q(
        POPCNT_5) );
    zdffqrb POPCNT_reg_4 ( .CK(CLK60M), .D(POPCNT1095_4), .R(STSRST_), .Q(
        POPCNT_4) );
    zdffqrb POPCNT_reg_3 ( .CK(CLK60M), .D(POPCNT1095_3), .R(STSRST_), .Q(
        POPCNT_3) );
    zdffqrb POPCNT_reg_2 ( .CK(CLK60M), .D(POPCNT1095_2), .R(STSRST_), .Q(
        POPCNT_2) );
    zdffqrb POPCNT_reg_1 ( .CK(CLK60M), .D(POPCNT1095_1), .R(STSRST_), .Q(
        POPCNT_1) );
    zdffqrb POPCNT_reg_0 ( .CK(CLK60M), .D(POPCNT1095_0), .R(STSRST_), .Q(
        POPCNT_0) );
    zivb U871 ( .A(POPCNT_0), .Y(POPCNT1087_0) );
    zdffqrb_ TX_HOSTDAT_reg_7 ( .CK(CLK60M), .D(TX_HOSTDAT1397_7), .R(TRST_), 
        .Q(TX_HOSTDAT_7) );
    zdffqrb_ TX_HOSTDAT_reg_6 ( .CK(CLK60M), .D(TX_HOSTDAT1397_6), .R(TRST_), 
        .Q(TX_HOSTDAT_6) );
    zdffqrb_ TX_HOSTDAT_reg_5 ( .CK(CLK60M), .D(TX_HOSTDAT1397_5), .R(TRST_), 
        .Q(TX_HOSTDAT_5) );
    zdffqrb_ TX_HOSTDAT_reg_4 ( .CK(CLK60M), .D(TX_HOSTDAT1397_4), .R(TRST_), 
        .Q(TX_HOSTDAT_4) );
    zdffqrb_ TX_HOSTDAT_reg_3 ( .CK(CLK60M), .D(TX_HOSTDAT1397_3), .R(TRST_), 
        .Q(TX_HOSTDAT_3) );
    zdffqrb_ TX_HOSTDAT_reg_2 ( .CK(CLK60M), .D(TX_HOSTDAT1397_2), .R(TRST_), 
        .Q(TX_HOSTDAT_2) );
    zdffqrb_ TX_HOSTDAT_reg_1 ( .CK(CLK60M), .D(TX_HOSTDAT1397_1), .R(TRST_), 
        .Q(TX_HOSTDAT_1) );
    zdffqsb EOPCNT_reg_0 ( .CK(CLK60M), .D(EOPCNT874_0), .S(TRST_), .Q(
        EOPCNT_0) );
    zdffqrb TXVALID_reg ( .CK(CLK60M), .D(TXVALID658), .R(TRST_), .Q(TXVALID)
         );
    zivb U872 ( .A(TXVALID), .Y(n2170) );
    zdffqrb TXSM_reg_6 ( .CK(CLK60M), .D(TXSM350_6), .R(TRST_), .Q(TXSM_6) );
    zivb U873 ( .A(TXSM_6), .Y(n2157) );
    zdffqrb PKTXEND_T_reg ( .CK(CLK60M), .D(n2252), .R(TRST_), .Q(PKTXEND_T)
         );
    zdffqrb_ TURNCNT_EN_reg ( .CK(CLK60M), .D(TURNCNT_EN488), .R(TRST_), .Q(
        TURNCNT_EN) );
    zdffqrb BYTECNT_reg_1 ( .CK(CLK60M), .D(BYTECNT836_1), .R(BYTECNTRST_), 
        .Q(BYTECNT_1) );
    zivb U874 ( .A(BYTECNT_1), .Y(n2076) );
    zdffqrb TXSM_reg_1 ( .CK(CLK60M), .D(TXSM350_1), .R(TRST_), .Q(TXSM_1) );
    zivb U875 ( .A(TXSM_1), .Y(n2151) );
    zdffqrb_ TXCRCEN_reg ( .CK(CLK60M), .D(val810_1), .R(TRST_), .Q(TXCRCEN)
         );
    zdffqsb TXSM_reg_0 ( .CK(CLK60M), .D(TXSM350_0), .S(TRST_), .Q(TXSM_0) );
    zivb U876 ( .A(TXSM_0), .Y(n2158) );
    zdffsb BYTECNT_reg_0 ( .CK(CLK60M), .D(BYTECNT836_0), .S(BYTECNTRST_), .Q(
        BYTECNT_0), .QN(n2074) );
    zdffqrb START_reg ( .CK(CLK60M), .D(START621), .R(TRST_), .Q(START) );
    zivb U877 ( .A(START), .Y(n2057) );
    zdffqrb PKTXEND_reg ( .CK(CLK60M), .D(n2250), .R(TRST_), .Q(PKTXEND) );
    zdffqrb TXRDY_reg ( .CK(CLK60M), .D(n1968), .R(TRST_), .Q(TXRDY) );
    zdffqrb SOF_DISCONN_P3_reg ( .CK(CLK60M), .D(n2248), .R(TRST_), .Q(
        SOF_DISCONN_P3) );
    zdffqrb PKTXEND_3T_reg ( .CK(CLK60M), .D(n2247), .R(TRST_), .Q(PKTXEND_3T)
         );
    zdffqrb SOF_DISCONN_P_reg ( .CK(CLK60M), .D(n2245), .R(TRST_), .Q(
        SOF_DISCONN_P) );
    zdffqrb TXCRC16_T_reg ( .CK(CLK60M), .D(USBPOP), .R(TRST_), .Q(TXCRC16_T)
         );
    zdffqrb_ TXCRCRST_reg ( .CK(CLK60M), .D(TXSM_0), .R(TRST_), .Q(TXCRCRST)
         );
    zdffqrb TEST_STATE_reg ( .CK(CLK60M), .D(TEST_STATE310), .R(TRST_), .Q(
        n1685) );
    zdffqrb PKTXEND_2T_reg ( .CK(CLK60M), .D(val1280_1), .R(TRST_), .Q(
        PKTXEND_2T) );
    zdffqrb SOF_DISCONN_T_reg ( .CK(CLK60M), .D(SOF_CHK_COND), .R(TRST_), .Q(
        SOF_DISCONN_T) );
    zdffrb BYTECNT_reg_2 ( .CK(CLK60M), .D(BYTECNT836_2), .R(BYTECNTRST_), .Q(
        BYTECNT_2), .QN(n2077) );
    zdffqrb SOF_DISCONN_P2_reg ( .CK(CLK60M), .D(n2243), .R(TRST_), .Q(
        SOF_DISCONN_P2) );
    zdffqrb PKTXEND_4T_reg ( .CK(CLK60M), .D(n1925), .R(TRST_), .Q(PKTXEND_4T)
         );
    zdffqrb EOPCNT_reg_4 ( .CK(CLK60M), .D(EOPCNT874_4), .R(TRST_), .Q(
        EOPCNT_4) );
    zivb U878 ( .A(EOPCNT_4), .Y(n1982) );
    zdffqrb TXSM_reg_2 ( .CK(CLK60M), .D(TXSM350_2), .R(TRST_), .Q(TXSM_2) );
    zivb U879 ( .A(TXSM_2), .Y(n2125) );
    zdffqrb TXSTART_T_reg ( .CK(CLK60M), .D(TXSTART_T584), .R(TRST_), .Q(
        TXSTART_T) );
    zivb U880 ( .A(TXSTART_T), .Y(n2059) );
    zdffqrb TEST_FLAG_reg ( .CK(CLK60M), .D(TEST_FLAG1306), .R(TRST_), .Q(
        TEST_FLAG) );
    zdffqrb TXSM_reg_3 ( .CK(CLK60M), .D(TXSM350_3), .R(TRST_), .Q(TXSM_3) );
    zivb U881 ( .A(TXSM_3), .Y(n1972) );
    zdffqrb TXCRC5_T_reg ( .CK(CLK60M), .D(TXCRC5_T732), .R(TRST_), .Q(
        TXCRC5_T) );
    zdffqrb TXSM_reg_4 ( .CK(CLK60M), .D(TXSM350_4), .R(TRST_), .Q(TXSM_4) );
    zivb U882 ( .A(TXSM_4), .Y(n2065) );
    znr2b U883 ( .A(TXSM_0), .B(n1932), .Y(n1925) );
    znr4b U884 ( .A(TXSM_4), .B(TXSM_1), .C(n2157), .D(n2156), .Y(n1926) );
    zan3b U885 ( .A(SPLIT), .B(n1934), .C(n2115), .Y(n1927) );
    znr2b U886 ( .A(n1960), .B(n2195), .Y(n1928) );
    znr2b U887 ( .A(SL_TXDATASEL[2]), .B(n1960), .Y(n1929) );
    zan3b U888 ( .A(n1934), .B(n1980), .C(n2115), .Y(n1930) );
    znr2b U889 ( .A(n2241), .B(n1935), .Y(n1931) );
    znr3b U890 ( .A(n2153), .B(n2200), .C(n2121), .Y(n1932) );
    znr4b U891 ( .A(TURN_CNT_1), .B(TURN_CNT_0), .C(TURN_CNT_2), .D(TURN_CNT_3
        ), .Y(n1933) );
    ziv11b U892 ( .A(n1990), .Y(n1934), .Z(n1935) );
    zivb U893 ( .A(TXCRCPHASE), .Y(n2067) );
    zdffqrb TXSM_reg_5 ( .CK(CLK60M), .D(TXSM350_5), .R(TRST_), .Q(TXCRCPHASE)
         );
    zdffrb EOPCNT_reg_3 ( .CK(CLK60M), .D(EOPCNT874_3), .R(TRST_), .QN(n1936)
         );
    zdffrb EOPCNT_reg_2 ( .CK(CLK60M), .D(EOPCNT874_2), .R(TRST_), .QN(n1937)
         );
    zdffrb EOPCNT_reg_1 ( .CK(CLK60M), .D(EOPCNT874_1), .R(TRST_), .Q(n2055), 
        .QN(n1938) );
    zor2b U894 ( .A(TXSM_2), .B(n2160), .Y(n2161) );
    zivb U895 ( .A(n2161), .Y(n2155) );
    zivb U896 ( .A(n2063), .Y(n2168) );
    znd2b U897 ( .A(n2235), .B(n1969), .Y(n2063) );
    zan2b U898 ( .A(n2050), .B(n1967), .Y(n1939) );
    znd2b U899 ( .A(n1975), .B(n1976), .Y(n2126) );
    zivb U900 ( .A(n2126), .Y(n2133) );
    znd3b U901 ( .A(n2067), .B(TXSM_3), .C(n2155), .Y(n2138) );
    zivb U902 ( .A(n2138), .Y(n2131) );
    zan2b U903 ( .A(n1955), .B(n2177), .Y(n1940) );
    zan2b U904 ( .A(n1955), .B(n2236), .Y(n1941) );
    zdffqrb_ TX_HOSTDAT_reg_0 ( .CK(CLK60M), .D(TX_HOSTDAT1397_0), .R(TRST_), 
        .Q(sub_551_carry_1) );
    zivb U905 ( .A(sub_551_carry_1), .Y(TX_HOSTDAT_N1348_0) );
    zivb U906 ( .A(n2115), .Y(n1942) );
    zan2b U907 ( .A(MACDATA_30), .B(n1942), .Y(n2113) );
    zan2b U908 ( .A(MACDATA_26), .B(n2241), .Y(n2109) );
    zan2b U909 ( .A(MACDATA_24), .B(n2241), .Y(n2107) );
    zan2b U910 ( .A(MACDATA_28), .B(n1942), .Y(n2111) );
    zao22b U911 ( .A(n1927), .B(CRC[3]), .C(MACDATA_22), .D(n1942), .Y(n2105)
         );
    zao22b U912 ( .A(ADRENDPS[17]), .B(n1927), .C(n1942), .D(MACDATA_17), .Y(
        n2100) );
    zao22b U913 ( .A(CRC[1]), .B(n1927), .C(MACDATA_20), .D(n1942), .Y(n2103)
         );
    zao22b U914 ( .A(ADRENDPS[18]), .B(n1927), .C(MACDATA_18), .D(n1942), .Y(
        n2101) );
    zan2b U915 ( .A(MACDATA_9), .B(n2241), .Y(n2139) );
    zmux21hb U916 ( .A(n2220), .B(MACDATA_2), .S(n2241), .Y(MACDATA388_2) );
    zmux21hb U917 ( .A(n2214), .B(MACDATA_4), .S(n2241), .Y(MACDATA388_4) );
    zmux21hb U918 ( .A(n2208), .B(MACDATA_6), .S(n2241), .Y(MACDATA388_6) );
    zor2b U919 ( .A(n2140), .B(n2171), .Y(n2237) );
    zmux21lb U920 ( .A(n2226), .B(MACDATA_0), .S(n2140), .Y(n2080) );
    zor2b U921 ( .A(n2140), .B(n2172), .Y(n2175) );
    zor2b U922 ( .A(n2056), .B(NXTISSYNC), .Y(n2115) );
    zivb U923 ( .A(n2115), .Y(n2140) );
    zdl1d U924 ( .A(n1963), .Y(n1943) );
    zdl1d U925 ( .A(n1966), .Y(n1944) );
    zxo2b U926 ( .A(POPCNT_5), .B(n1953), .Y(n2044) );
    zbfp U927 ( .A(MAXLEN[5]), .Y(n1953) );
    znr5d U928 ( .A(n2033), .B(n1917), .C(n1920), .D(n1923), .E(n1924), .Y(
        n1945) );
    zbfh U929 ( .A(MAXLEN[4]), .Y(n1946) );
    zivb U930 ( .A(n1949), .Y(n2201) );
    zdl1d U931 ( .A(MAXLEN[6]), .Y(n1965) );
    zdl1d U932 ( .A(n2016), .Y(n1947) );
    znr2d U933 ( .A(n1958), .B(n1948), .Y(n1954) );
    zivl U934 ( .A(n2020), .Y(n1948) );
    zivb U935 ( .A(n1958), .Y(n1964) );
    znd2b U936 ( .A(n1945), .B(n2018), .Y(n1958) );
    zdl1d U937 ( .A(n2023), .Y(n1949) );
    zbfh U938 ( .A(MAXLEN[1]), .Y(n1950) );
    zbfh U939 ( .A(MAXLEN[10]), .Y(n1952) );
    zan2b U940 ( .A(n1964), .B(n2020), .Y(n1955) );
    zmux21lb U941 ( .A(n1961), .B(n2125), .S(n2168), .Y(TXSM350_2) );
    zor2b U942 ( .A(TXSM_2), .B(n1961), .Y(n2178) );
    zbfh U943 ( .A(MAXLEN[8]), .Y(n1956) );
    znr6d U944 ( .A(n2026), .B(n2013), .C(n2025), .D(n2029), .E(n2027), .F(
        n2028), .Y(n1957) );
    znr2b U945 ( .A(n1955), .B(n2012), .Y(n1988) );
    znd2b U946 ( .A(n2115), .B(n1955), .Y(n2176) );
    zaoi21b U947 ( .A(n1955), .B(n1983), .C(n1984), .Y(n2068) );
    zao21b U948 ( .A(SL_TXDATASEL[1]), .B(USBPOP), .C(TXSTART), .Y(n2070) );
    zmux21hb U949 ( .A(POPCNT_0), .B(POPCNT1087_0), .S(USBPOP), .Y(
        POPCNT1095_0) );
    zmux21hb U950 ( .A(POPCNT_1), .B(POPCNT1087_1), .S(USBPOP), .Y(
        POPCNT1095_1) );
    zmux21hb U951 ( .A(POPCNT_10), .B(POPCNT1087_10), .S(USBPOP), .Y(
        POPCNT1095_10) );
    zmux21hb U952 ( .A(POPCNT_2), .B(POPCNT1087_2), .S(USBPOP), .Y(
        POPCNT1095_2) );
    zmux21hb U953 ( .A(POPCNT_3), .B(POPCNT1087_3), .S(USBPOP), .Y(
        POPCNT1095_3) );
    zmux21hb U954 ( .A(POPCNT_4), .B(POPCNT1087_4), .S(USBPOP), .Y(
        POPCNT1095_4) );
    zmux21hb U955 ( .A(POPCNT_5), .B(POPCNT1087_5), .S(USBPOP), .Y(
        POPCNT1095_5) );
    zmux21hb U956 ( .A(POPCNT_6), .B(POPCNT1087_6), .S(USBPOP), .Y(
        POPCNT1095_6) );
    zmux21hb U957 ( .A(POPCNT_7), .B(POPCNT1087_7), .S(USBPOP), .Y(
        POPCNT1095_7) );
    zmux21hb U958 ( .A(POPCNT_8), .B(POPCNT1087_8), .S(USBPOP), .Y(
        POPCNT1095_8) );
    zmux21hb U959 ( .A(POPCNT_9), .B(POPCNT1087_9), .S(USBPOP), .Y(
        POPCNT1095_9) );
    zor2b U960 ( .A(TXSTART), .B(USBPOP), .Y(n2165) );
    zdffrb_ USBPOP_reg ( .CK(CLK60M), .D(USBPOP1137), .R(STSRST_), .Q(USBPOP), 
        .QN(n1960) );
    zdl1d U961 ( .A(n2169), .Y(n1961) );
    zbfh U962 ( .A(MAXLEN[0]), .Y(n1962) );
    zbfh U963 ( .A(MAXLEN[9]), .Y(n1966) );
    znd2b U964 ( .A(n1964), .B(n2020), .Y(n1967) );
    ziv22b U965 ( .A(TXREADY), .Y1(n1969), .Y2(n1968) );
    zind2d U966 ( .A(n2154), .B(n1973), .Y(n2156) );
    znd2d U967 ( .A(n2063), .B(n1977), .Y(n2064) );
    zcx1d U968 ( .A(n1978), .B(n1979), .C(n2063), .D(n1972), .Y(TXSM350_3) );
    znd2d U969 ( .A(n2056), .B(n1967), .Y(n2075) );
    zcxi2d U970 ( .A(n2120), .B(n1938), .C(EOPCNT_0), .D(n2117), .Y(
        EOPCNT874_1) );
    zcxi2d U971 ( .A(n2120), .B(n1937), .C(n2055), .D(n2117), .Y(EOPCNT874_2)
         );
    zoai22d U972 ( .A(n2120), .B(n1936), .C(n1981), .D(n1937), .Y(EOPCNT874_3)
         );
    zoai22d U973 ( .A(n2120), .B(n1982), .C(n1981), .D(n1936), .Y(EOPCNT874_4)
         );
    zaoi21d U974 ( .A(n2201), .B(n2133), .C(n1988), .Y(n2066) );
    znd6d U975 ( .A(n2054), .B(n1990), .C(n1967), .D(n2235), .E(n2171), .F(
        n2178), .Y(n2172) );
    zoai21d U976 ( .A(n2007), .B(n2008), .C(n1977), .Y(n2169) );
    zaoi21d U977 ( .A(n2169), .B(n2054), .C(n2009), .Y(USBPOP1137) );
    znr4d U978 ( .A(n1954), .B(n2010), .C(n2126), .D(HANDSHK), .Y(n2007) );
    zinr2b U979 ( .A(TX_PID[0]), .B(n2178), .Y(n1992) );
    zxo2d U980 ( .A(TXBCNT[0]), .B(n1962), .Y(n2013) );
    zivh U981 ( .A(DATPKT), .Y(n2015) );
    znd2d U982 ( .A(n1957), .B(n2017), .Y(n2016) );
    znd2d U983 ( .A(TOKEN), .B(TXSM_2), .Y(n1990) );
    znd2d U984 ( .A(DIS_STUFF), .B(n1968), .Y(n1981) );
    znd2d U985 ( .A(n1947), .B(n2019), .Y(n1989) );
    znd2d U986 ( .A(n2016), .B(n2024), .Y(n2023) );
    zxo2d U987 ( .A(TXBCNT[9]), .B(n1966), .Y(n2025) );
    zxo2d U988 ( .A(TXBCNT[6]), .B(MAXLEN[6]), .Y(n2026) );
    zxo2d U989 ( .A(n1952), .B(TXBCNT[10]), .Y(n2027) );
    zxo2d U990 ( .A(n1951), .B(TXBCNT[2]), .Y(n2028) );
    zxo2d U991 ( .A(n1950), .B(TXBCNT[1]), .Y(n2029) );
    zxo2d U992 ( .A(TXBCNT[3]), .B(n1963), .Y(n2030) );
    zxo2d U993 ( .A(n1953), .B(TXBCNT[5]), .Y(n2031) );
    zxo2d U994 ( .A(TXBCNT[8]), .B(n1956), .Y(n2032) );
    zxo2d U995 ( .A(TXBCNT[7]), .B(MAXLEN[7]), .Y(n2033) );
    zxo2d U996 ( .A(TXBCNT[4]), .B(n1946), .Y(n2034) );
    zxo2d U997 ( .A(n1944), .B(POPCNT_9), .Y(n2035) );
    zxo2d U998 ( .A(POPCNT_3), .B(n1943), .Y(n2037) );
    zxo2d U999 ( .A(POPCNT_10), .B(n1952), .Y(n2040) );
    zxo2d U1000 ( .A(POPCNT_8), .B(n1956), .Y(n2041) );
    zxo2d U1001 ( .A(POPCNT_1), .B(n1950), .Y(n2042) );
    zxo2d U1002 ( .A(POPCNT_2), .B(n1951), .Y(n2043) );
    znr6d U1003 ( .A(n1918), .B(n2026), .C(n1921), .D(n2029), .E(n1919), .F(
        n1922), .Y(n2018) );
    znr5d U1004 ( .A(n2033), .B(n2034), .C(n2032), .D(n2030), .E(n2031), .Y(
        n2017) );
    znr6d U1005 ( .A(n2014), .B(n2036), .C(n2035), .D(n2039), .E(n2037), .F(
        n2038), .Y(n2045) );
    znr5d U1006 ( .A(n2043), .B(n2044), .C(n2042), .D(n2040), .E(n2041), .Y(
        n2046) );
    znr3d U1007 ( .A(n1969), .B(n2015), .C(n2047), .Y(n2024) );
    znd2d U1008 ( .A(n2023), .B(n1990), .Y(n2010) );
    zinr2b U1009 ( .A(n2158), .B(TXSM_2), .Y(n1973) );
    zcxi2d U1010 ( .A(n1968), .B(n2126), .C(n2048), .D(BYTECNT_3), .Y(n2008)
         );
    znr2d U1011 ( .A(n2015), .B(n2047), .Y(n2019) );
    zcx3d U1012 ( .A(n2046), .B(n2045), .C(n2049), .D(TXRDY), .Y(n2009) );
    znd2d U1013 ( .A(DATPKT), .B(TXSM_2), .Y(n2051) );
    znd2d U1014 ( .A(n2065), .B(n2051), .Y(n2020) );
    zor2d U1015 ( .A(TXSM_4), .B(TXSM_2), .Y(n2052) );
    zivf U1016 ( .A(n2052), .Y(n2047) );
    zcxi2d U1017 ( .A(n2126), .B(n1990), .C(n2053), .D(n2131), .Y(n1978) );
    zind2d U1018 ( .A(n2054), .B(HOSTTMP_1), .Y(n2006) );
    zind2d U1019 ( .A(n2054), .B(HOSTTMP_2), .Y(n2004) );
    zind2d U1020 ( .A(n2054), .B(HOSTTMP_3), .Y(n2002) );
    zind2d U1021 ( .A(n2054), .B(HOSTTMP_4), .Y(n2000) );
    zind2d U1022 ( .A(n2054), .B(HOSTTMP_5), .Y(n1998) );
    zind2d U1023 ( .A(n2054), .B(HOSTTMP_6), .Y(n1996) );
    zind2d U1024 ( .A(n2054), .B(HOSTTMP_7), .Y(n1994) );
    zbfp U1025 ( .A(n1989), .Y(n2054) );
    zdffqrb BYTECNT_reg_3 ( .CK(CLK60M), .D(BYTECNT836_3), .R(BYTECNTRST_), 
        .Q(BYTECNT_3) );
    zdffqrd TXBCNT_reg_5 ( .CK(CLK60M), .D(TXBCNT446_5), .R(TXBCNTRST_), .Q(
        TXBCNT[5]) );
    zdffqrd TXBCNT_reg_3 ( .CK(CLK60M), .D(TXBCNT446_3), .R(TXBCNTRST_), .Q(
        TXBCNT[3]) );
    zhadrd add_272_U1_1_5 ( .A(TXBCNT[5]), .B(add_272_carry_5), .CO(
        add_272_carry_6), .S(TXBCNT438_5) );
    zhadrd add_272_U1_1_3 ( .A(TXBCNT[3]), .B(add_272_carry_3), .CO(
        add_272_carry_4), .S(TXBCNT438_3) );
    zor3b U1026 ( .A(TXSM_6), .B(n1685), .C(SL_FORCE_STUFF), .Y(DIS_STUFF) );
    zor4b U1027 ( .A(TEST_K), .B(n1685), .C(TEST_EYE), .D(TEST_J), .Y(
        TEST_STATE310) );
    zoa21d U1029 ( .A(TEST_J), .B(TEST_FLAG), .C(n_2889), .Y(n_2892) );
    zor3b U1030 ( .A(START), .B(n1685), .C(n1932), .Y(TXVALID658) );
    zao222b U1031 ( .A(TXCRCDAT[7]), .B(n1960), .C(HOSTDAT[7]), .D(n1929), .E(
        n1928), .F(TX_HOSTDAT_7), .Y(HOSTD978_7) );
    zao222b U1032 ( .A(TXCRCDAT[6]), .B(n1960), .C(HOSTDAT[6]), .D(n1929), .E(
        n1928), .F(TX_HOSTDAT_6), .Y(HOSTD978_6) );
    zao222b U1033 ( .A(TXCRCDAT[5]), .B(n1960), .C(HOSTDAT[5]), .D(n1929), .E(
        n1928), .F(TX_HOSTDAT_5), .Y(HOSTD978_5) );
    zao222b U1034 ( .A(TXCRCDAT[4]), .B(n1960), .C(HOSTDAT[4]), .D(n1929), .E(
        n1928), .F(TX_HOSTDAT_4), .Y(HOSTD978_4) );
    zao222b U1035 ( .A(TXCRCDAT[3]), .B(n1960), .C(HOSTDAT[3]), .D(n1929), .E(
        n1928), .F(TX_HOSTDAT_3), .Y(HOSTD978_3) );
    zao222b U1036 ( .A(TXCRCDAT[2]), .B(n1960), .C(HOSTDAT[2]), .D(n1929), .E(
        n1928), .F(TX_HOSTDAT_2), .Y(HOSTD978_2) );
    zao222b U1037 ( .A(TXCRCDAT[1]), .B(n1960), .C(HOSTDAT[1]), .D(n1929), .E(
        n1928), .F(TX_HOSTDAT_1), .Y(HOSTD978_1) );
    zao222b U1038 ( .A(TXCRCDAT[0]), .B(n1960), .C(HOSTDAT[0]), .D(n1929), .E(
        n1928), .F(sub_551_carry_1), .Y(HOSTD978_0) );
    zoa21d U1039 ( .A(n2062), .B(DIS_NARROW_SOF), .C(SOF_DISCONN_P), .Y(
        SOF_DISCONN) );
    zoai22d U1040 ( .A(n2065), .B(n2063), .C(n2066), .D(n2064), .Y(TXSM350_4)
         );
    zoai22d U1041 ( .A(n2067), .B(n2063), .C(n2068), .D(n2064), .Y(TXSM350_5)
         );
    zoai211d U1042 ( .A(n2073), .B(n2074), .C(TXVALID), .D(n1939), .Y(
        BYTECNT836_0) );
    zoai22d U1043 ( .A(n2075), .B(n2074), .C(n2076), .D(n2073), .Y(
        BYTECNT836_1) );
    zoai22d U1044 ( .A(n2076), .B(n2075), .C(n2077), .D(n2073), .Y(
        BYTECNT836_2) );
    zoai22d U1045 ( .A(n2077), .B(n2075), .C(n2078), .D(n2073), .Y(
        BYTECNT836_3) );
    zao211b U1046 ( .A(MACDATA_16), .B(n2079), .C(n2082), .D(n2083), .Y(
        MACDATA388_8) );
    zao211b U1047 ( .A(MACDATA_17), .B(n2240), .C(n2084), .D(n2085), .Y(
        MACDATA388_9) );
    zao211b U1048 ( .A(MACDATA_18), .B(n2079), .C(n2086), .D(n2087), .Y(
        MACDATA388_10) );
    zao211b U1049 ( .A(MACDATA_19), .B(n2240), .C(n2088), .D(n2089), .Y(
        MACDATA388_11) );
    zao211b U1050 ( .A(MACDATA_20), .B(n2079), .C(n2090), .D(n2091), .Y(
        MACDATA388_12) );
    zao211b U1051 ( .A(MACDATA_21), .B(n2240), .C(n2092), .D(n2093), .Y(
        MACDATA388_13) );
    zao211b U1052 ( .A(MACDATA_22), .B(n2079), .C(n2094), .D(n2095), .Y(
        MACDATA388_14) );
    zao211b U1053 ( .A(MACDATA_23), .B(n2240), .C(n2096), .D(n2097), .Y(
        MACDATA388_15) );
    zao211b U1054 ( .A(MACDATA_24), .B(n2079), .C(n2098), .D(n2242), .Y(
        MACDATA388_16) );
    zao211b U1055 ( .A(MACDATA_25), .B(n2240), .C(n2100), .D(n2099), .Y(
        MACDATA388_17) );
    zao211b U1056 ( .A(MACDATA_26), .B(n2079), .C(n2101), .D(n2242), .Y(
        MACDATA388_18) );
    zao211b U1057 ( .A(MACDATA_27), .B(n2240), .C(n2102), .D(n2099), .Y(
        MACDATA388_19) );
    zao211b U1058 ( .A(MACDATA_28), .B(n2079), .C(n2103), .D(n2242), .Y(
        MACDATA388_20) );
    zao211b U1059 ( .A(MACDATA_29), .B(n2240), .C(n2104), .D(n2099), .Y(
        MACDATA388_21) );
    zao211b U1060 ( .A(MACDATA_30), .B(n2079), .C(n2105), .D(n2242), .Y(
        MACDATA388_22) );
    zao211b U1061 ( .A(MACDATA_31), .B(n2240), .C(n2106), .D(n2099), .Y(
        MACDATA388_23) );
    zao211b U1062 ( .A(MACDATA_32), .B(n2079), .C(n2099), .D(n2107), .Y(
        MACDATA388_24) );
    zao211b U1063 ( .A(MACDATA_33), .B(n2240), .C(n2242), .D(n2108), .Y(
        MACDATA388_25) );
    zao211b U1064 ( .A(MACDATA_34), .B(n2079), .C(n2099), .D(n2109), .Y(
        MACDATA388_26) );
    zao211b U1065 ( .A(MACDATA_35), .B(n2240), .C(n2242), .D(n2110), .Y(
        MACDATA388_27) );
    zao211b U1066 ( .A(MACDATA_36), .B(n2079), .C(n2099), .D(n2111), .Y(
        MACDATA388_28) );
    zao211b U1067 ( .A(MACDATA_37), .B(n2240), .C(n2099), .D(n2112), .Y(
        MACDATA388_29) );
    zao211b U1068 ( .A(MACDATA_38), .B(n2079), .C(n2242), .D(n2113), .Y(
        MACDATA388_30) );
    zoa21d U1069 ( .A(TURNCNT_EN), .B(PKTXEND), .C(n2116), .Y(TURNCNT_EN488)
         );
    zao211b U1070 ( .A(EOPCNT_4), .B(n2117), .C(n2118), .D(n2119), .Y(
        EOPCNT874_0) );
    zoa21d U1071 ( .A(n2118), .B(n2128), .C(SOF_DISCONN_CHK), .Y(n2058) );
    zan2d U1072 ( .A(EOPCNT_0), .B(n2150), .Y(n2119) );
    zoai21d U1073 ( .A(n2151), .B(n2063), .C(n2152), .Y(TXSM350_1) );
    zor4b U1074 ( .A(TXSM_2), .B(n2158), .C(n2154), .D(n2159), .Y(n2136) );
    zor3b U1075 ( .A(n1960), .B(n2162), .C(SL_TXDATASEL[1]), .Y(n2163) );
    zor3b U1076 ( .A(n1960), .B(SL_TXDATASEL[0]), .C(SL_TXDATASEL[1]), .Y(
        n2164) );
    zor3b U1077 ( .A(n2170), .B(n1968), .C(n1955), .Y(n2073) );
    zmux21ld U1078 ( .A(n2167), .B(n2157), .S(n2168), .Y(TXSM350_6) );
    zmux21ld U1079 ( .A(n1932), .B(n2158), .S(n2168), .Y(TXSM350_0) );
    zmux21hd U1080 ( .A(TXBCNT[9]), .B(TXBCNT438_9), .S(n2201), .Y(TXBCNT446_9
        ) );
    zmux21hd U1081 ( .A(TXBCNT[8]), .B(TXBCNT438_8), .S(n2201), .Y(TXBCNT446_8
        ) );
    zmux21hd U1082 ( .A(TXBCNT[7]), .B(TXBCNT438_7), .S(n2201), .Y(TXBCNT446_7
        ) );
    zmux21hd U1083 ( .A(TXBCNT[6]), .B(TXBCNT438_6), .S(n2201), .Y(TXBCNT446_6
        ) );
    zmux21hd U1084 ( .A(TXBCNT[5]), .B(TXBCNT438_5), .S(n2201), .Y(TXBCNT446_5
        ) );
    zmux21hd U1085 ( .A(TXBCNT[4]), .B(TXBCNT438_4), .S(n2201), .Y(TXBCNT446_4
        ) );
    zmux21hd U1086 ( .A(TXBCNT[3]), .B(TXBCNT438_3), .S(n2201), .Y(TXBCNT446_3
        ) );
    zmux21hd U1087 ( .A(TXBCNT[2]), .B(TXBCNT438_2), .S(n2201), .Y(TXBCNT446_2
        ) );
    zmux21hd U1088 ( .A(TXBCNT[10]), .B(TXBCNT438_10), .S(n2201), .Y(
        TXBCNT446_10) );
    zmux21hd U1089 ( .A(TXBCNT[1]), .B(TXBCNT438_1), .S(n2201), .Y(TXBCNT446_1
        ) );
    zmux21hd U1090 ( .A(TXBCNT[0]), .B(TXBCNT438_0), .S(n2201), .Y(TXBCNT446_0
        ) );
    zao211b U1091 ( .A(MACDATA_15), .B(n2205), .C(n2206), .D(n2207), .Y(n2204)
         );
    zao211b U1092 ( .A(MACDATA_14), .B(n2205), .C(n2209), .D(n2210), .Y(n2208)
         );
    zao211b U1093 ( .A(MACDATA_13), .B(n2205), .C(n2212), .D(n2213), .Y(n2211)
         );
    zao211b U1094 ( .A(MACDATA_12), .B(n2205), .C(n2215), .D(n2216), .Y(n2214)
         );
    zao211b U1095 ( .A(MACDATA_11), .B(n2205), .C(n2218), .D(n2219), .Y(n2217)
         );
    zao211b U1096 ( .A(MACDATA_10), .B(n2205), .C(n2221), .D(n2222), .Y(n2220)
         );
    zao211b U1097 ( .A(MACDATA_9), .B(n2205), .C(n2224), .D(n2225), .Y(n2223)
         );
    zao211b U1098 ( .A(TXSM_0), .B(n2159), .C(n2166), .D(n2123), .Y(n2227) );
    zao222b U1099 ( .A(TXSM_4), .B(TXSM_6), .C(TXCRCPHASE), .D(TXSM_3), .E(
        n2229), .F(n2057), .Y(n2228) );
    zao211b U1100 ( .A(TXSM_2), .B(n2160), .C(n2227), .D(n2228), .Y(n2200) );
    zao211b U1101 ( .A(ADRENDPS[9]), .B(n1931), .C(n2242), .D(n2139), .Y(n2084
        ) );
    zao211b U1102 ( .A(ADRENDPS[8]), .B(n1931), .C(n2099), .D(n2141), .Y(n2082
        ) );
    zao211b U1103 ( .A(n2174), .B(TX_PID[7]), .C(n2173), .D(n2142), .Y(n2207)
         );
    zao211b U1104 ( .A(TX_PID[6]), .B(n2174), .C(n2173), .D(n2143), .Y(n2210)
         );
    zao211b U1105 ( .A(TX_PID[5]), .B(n2174), .C(n2173), .D(n2144), .Y(n2213)
         );
    zao211b U1106 ( .A(TX_PID[4]), .B(n2174), .C(n2173), .D(n2145), .Y(n2216)
         );
    zao211b U1107 ( .A(MACDATA_31), .B(n1942), .C(NXTISSYNC), .D(n2242), .Y(
        n2114) );
    zao211b U1108 ( .A(TX_PID[3]), .B(n2174), .C(n2173), .D(n2146), .Y(n2219)
         );
    zao211b U1109 ( .A(TX_PID[2]), .B(n2174), .C(n2173), .D(n2147), .Y(n2222)
         );
    zao211b U1110 ( .A(MACDATA_15), .B(n1942), .C(n2099), .D(n2230), .Y(n2097)
         );
    zao211b U1111 ( .A(MACDATA_14), .B(n2241), .C(n2242), .D(n2231), .Y(n2095)
         );
    zao211b U1112 ( .A(MACDATA_13), .B(n2241), .C(n2099), .D(n2232), .Y(n2093)
         );
    zao211b U1113 ( .A(MACDATA_12), .B(n1942), .C(n2242), .D(n2233), .Y(n2091)
         );
    zao211b U1114 ( .A(MACDATA_11), .B(n2241), .C(n2099), .D(n2234), .Y(n2089)
         );
    zao211b U1115 ( .A(ADRENDPS[10]), .B(n1931), .C(n2242), .D(n2148), .Y(
        n2086) );
    zao211b U1116 ( .A(TX_PID[1]), .B(n2174), .C(n2173), .D(n2149), .Y(n2225)
         );
    zao211b U1117 ( .A(BYTECNT_2), .B(SPLIT), .C(BYTECNT_0), .D(BYTECNT_1), 
        .Y(n2061) );
    zor4b U1118 ( .A(n2198), .B(n2199), .C(n2196), .D(n2197), .Y(n2116) );
    zor2d S_238 ( .A(n_4084), .B(ATPG_ENI), .Y(BYTECNTRST_) );
    zan2d S_237 ( .A(STSRST_), .B(n_4083), .Y(n_4084) );
    zan2d S_162 ( .A(STSRST_), .B(TXVALID), .Y(n_3829) );
    zor2d S_163 ( .A(n_3829), .B(ATPG_ENI), .Y(TXBCNTRST_) );
    zao21b U1119 ( .A(n1685), .B(n2056), .C(TEST_FLAG), .Y(TEST_FLAG1306) );
    zbfb U1120 ( .A(SOF_DISCONN_P), .Y(n2243) );
    zivb U1121 ( .A(SOF_DISCONN_T), .Y(n2244) );
    zivb U1122 ( .A(n2244), .Y(n2245) );
    zivb U1123 ( .A(PKTXEND_4T), .Y(n2246) );
    zivb U1124 ( .A(n2246), .Y(n2247) );
    zbfb U1125 ( .A(SOF_DISCONN_P2), .Y(n2248) );
    zivb U1126 ( .A(PKTXEND_T), .Y(n2249) );
    zivb U1127 ( .A(n2249), .Y(n2250) );
    zivb U1128 ( .A(PKTXEND_2T), .Y(n2251) );
    zivb U1129 ( .A(n2251), .Y(n2252) );
    zbfb U1130 ( .A(HOSTTMP1039_1), .Y(n2253) );
    zbfb U1131 ( .A(HOSTTMP1039_2), .Y(n2254) );
    zbfb U1132 ( .A(HOSTTMP1039_3), .Y(n2255) );
    zbfb U1133 ( .A(HOSTTMP1039_4), .Y(n2256) );
    zbfb U1134 ( .A(HOSTTMP1039_5), .Y(n2257) );
    zbfb U1135 ( .A(HOSTTMP1039_6), .Y(n2258) );
    zbfb U1136 ( .A(HOSTTMP1039_7), .Y(n2259) );
endmodule


module HS_RXCTL ( DATA_RX, RXACTIVE, RXVALID, CLK60M, ASKREPLY, TRST_, STSRST_, 
    USBDAT, PIDERR, RXPID, RXDATA, RXHAND, RXSTUFFERR, LATCHDAT, RXCRCEN, 
    RXCRCRST, RXCRCDAT, LATCHPID, CRCHK, PKRVEND, RXEOPERR, DISCHKEOPERR, 
    PHYERR, CRCERR, NORMPKT, EOF2, TMOUT, MAXLEN, BABBLE, RXBCNT, RXDATA0, 
    RXDATA1, RXDATA2, RXMDATA, DAT0, DAT1, DAT2, DATM, ISO, RXACK, TOGMATCH, 
    SPD, RXTOKENPHASE, DATAIN, RXSOF, RXTOKEN, RXADDRF, MAC_SLAVE_ACT, 
    SL_TOGMATCH, EXEITD, LATCHADDR, EN_CHKTOGCRC, EN_REF_RVLD, RVLD );
input  [7:0] DATA_RX;
output [7:0] USBDAT;
output [7:0] RXPID;
output [7:0] RXCRCDAT;
output [23:0] RXADDRF;
input  [10:0] MAXLEN;
output [10:0] RXBCNT;
input  RXACTIVE, RXVALID, CLK60M, ASKREPLY, TRST_, STSRST_, PIDERR, RXDATA, 
    RXHAND, RXSTUFFERR, RXEOPERR, DISCHKEOPERR, CRCERR, EOF2, TMOUT, RXDATA0, 
    RXDATA1, RXDATA2, RXMDATA, DAT0, DAT1, DAT2, DATM, ISO, RXACK, 
    RXTOKENPHASE, DATAIN, RXSOF, RXTOKEN, MAC_SLAVE_ACT, SL_TOGMATCH, EXEITD, 
    EN_CHKTOGCRC, EN_REF_RVLD, RVLD;
output LATCHDAT, RXCRCEN, RXCRCRST, LATCHPID, CRCHK, PKRVEND, PHYERR, NORMPKT, 
    BABBLE, TOGMATCH, SPD, LATCHADDR;
    wire RXACTIVE_FLAG, HOLD_14, RXBCNT981_2, RXVALID_L2H, RXPID535_0, 
        RXBCNT989_3, SPAREO6, n_2676, RXSM_0, ADDSEL1101_0, SPAREO0_, 
        PHYERR291, n_2277, SPAREO8, RVLD_SYNC, n_2678, n_2265, RXSTART, 
        LATCHDAT_P, RXBCNT989_4, SPAREO1, EN_LATCHDAT, RXBCNT981_5, HOLD_13, 
        RXPID535_7, n_1864, CRCEN_T624, RXSM457_0, SPAREO9, ADDSEL1101_1, 
        n_2670, RXSM_1, RXVALID_SYNC_T, HOLD_12, RXBCNT981_4, RXVALID_SYNC_2T, 
        RXPID535_6, RXSM457_1, RXBCNT989_5, SPAREO0, n_2263, RXBCNT989_2, 
        SPAREO7, HOLD_15, RXBCNT981_3, NXTISADR, LATCHDAT783, n_2680, n_1862, 
        RXPID535_1, n_1870, PKRVEND_T, RXBCNT989_10, n_2271, RXPID535_3, 
        n_1860, RXSM457_4, RXBCNT981_1, RXSTART587, SPAREO5, RXBCNT989_0, 
        val832_1, RXBCNT981_10, CRCEN_T, RXBCNT981_8, RXBCNT989_9, n_2273, 
        RXSM_4, RXSM_3, n_1872, n_2672, RXVALID_L2H736, SPAREO2, RXBCNT989_7, 
        RXSM457_3, RXPID535_4, HOLD_8, RXBCNT981_6, HOLD_10, n_2668, n_2275, 
        RXSM_2, ADDSEL1101_2, BABBLE1031, n_1874, RXSM457_2, n_1866, 
        RXPID535_5, HOLD_11, HOLD_9, RXBCNT981_7, SPAREO3, RXBCNT989_6, 
        SPAREO1_, n_2267, RXACTIVE_SYNC, n_2666, SPAREO4, RXBCNT989_1, 
        RXPID535_2, RXBCNT981_0, n_2269, n_2674, RXBCNT989_8, n_1868, 
        RXBCNT981_9, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
        n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
        n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
        n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
        n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
        n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
        n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
        n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
        n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
        add_377_carry_8, add_377_carry_6, add_377_carry_7, add_377_carry_9, 
        add_377_carry_2, add_377_carry_5, add_377_carry_10, add_377_carry_4, 
        add_377_carry_3, n1540, n1541, n1542, n1543, n1544, n1545, n1546, 
        n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, 
        n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, 
        n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, 
        n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, 
        n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, 
        n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, 
        n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, 
        n1617, n1618, n1619, n1620, n1621, n1622;
    zdffrb SPARE660 ( .CK(CLK60M), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE669 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb SPARE667 ( .A(SPAREO4), .Y(SPAREO5) );
    znr3b SPARE666 ( .A(SPAREO2), .B(n1536), .C(SPAREO0_), .Y(SPAREO4) );
    zdffrb SPARE661 ( .CK(CLK60M), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE668 ( .A(SPAREO5), .Y(SPAREO6) );
    zaoi211b SPARE663 ( .A(SPAREO4), .B(n1457), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zoai21b SPARE664 ( .A(SPAREO0), .B(SPAREO8), .C(EN_LATCHDAT), .Y(SPAREO9)
         );
    zoai21b SPARE665 ( .A(SPAREO1), .B(NXTISADR), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE662 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zan2b U458 ( .A(n1543), .B(n1549), .Y(NXTISADR) );
    znr6b U459 ( .A(RXBCNT[1]), .B(RXBCNT[9]), .C(RXBCNT[2]), .D(RXBCNT[4]), 
        .E(RXBCNT[5]), .F(RXBCNT[3]), .Y(n1503) );
    znr4b U460 ( .A(n1483), .B(RXBCNT[7]), .C(RXBCNT[8]), .D(RXBCNT[6]), .Y(
        n1502) );
    znd2b U461 ( .A(MAXLEN[0]), .B(RXBCNT981_0), .Y(n1508) );
    znd2b U462 ( .A(MAXLEN[2]), .B(n1478), .Y(n1510) );
    znd2b U463 ( .A(RXBCNT[2]), .B(n1489), .Y(n1524) );
    zivc U464 ( .A(MAXLEN[2]), .Y(n1489) );
    znd2b U465 ( .A(n1458), .B(n1483), .Y(n1518) );
    znd2b U466 ( .A(RXBCNT[0]), .B(n1482), .Y(n1517) );
    zivc U467 ( .A(MAXLEN[0]), .Y(n1482) );
    znd2b U468 ( .A(RXBCNT[7]), .B(n1484), .Y(n1516) );
    znd2b U469 ( .A(n1595), .B(n1461), .Y(n1469) );
    zor2b U470 ( .A(RXACTIVE_SYNC), .B(n1547), .Y(n1595) );
    zan3b U471 ( .A(n1568), .B(n1569), .C(n1570), .Y(n1567) );
    zivb U472 ( .A(RXTOKEN), .Y(n1579) );
    zan3b U473 ( .A(RXSM_0), .B(n1549), .C(n1452), .Y(n1566) );
    zor2b U474 ( .A(RXSTART), .B(RXACTIVE_SYNC), .Y(n1586) );
    zan2b U475 ( .A(n1584), .B(RXVALID), .Y(n1493) );
    znd2b U476 ( .A(RXDATA), .B(n1453), .Y(n1463) );
    znd2b U477 ( .A(RXACTIVE_SYNC), .B(n1587), .Y(n1462) );
    zivb U478 ( .A(n1585), .Y(n1587) );
    znd2b U479 ( .A(n1534), .B(n1535), .Y(n1466) );
    zivh U480 ( .A(EN_LATCHDAT), .Y(n1532) );
    zivb U481 ( .A(n1576), .Y(n1568) );
    zor2b U482 ( .A(n1578), .B(n1454), .Y(n1577) );
    zivb U483 ( .A(n1586), .Y(n1578) );
    znr2b U484 ( .A(n1582), .B(n1571), .Y(n1530) );
    znd2b U485 ( .A(n1573), .B(n1533), .Y(n1531) );
    zivb U486 ( .A(RXACK), .Y(n1533) );
    znr4b U487 ( .A(n1515), .B(n1519), .C(n1523), .D(n1527), .Y(n1496) );
    znd3b U488 ( .A(n1516), .B(n1517), .C(n1518), .Y(n1515) );
    znd3b U489 ( .A(n1520), .B(n1521), .C(n1522), .Y(n1519) );
    znd3b U490 ( .A(n1524), .B(n1525), .C(n1526), .Y(n1523) );
    znd2b U491 ( .A(n1528), .B(n1529), .Y(n1527) );
    zivb U492 ( .A(n1575), .Y(n1464) );
    zmux21hb U493 ( .A(RXBCNT[0]), .B(RXBCNT981_0), .S(LATCHDAT), .Y(
        RXBCNT989_0) );
    zao22b U494 ( .A(n1561), .B(n1544), .C(n1562), .D(RXSM_2), .Y(RXSM457_2)
         );
    zao21b U495 ( .A(n1456), .B(n1561), .C(n1468), .Y(RXSM457_1) );
    znr2b U496 ( .A(n1559), .B(n1560), .Y(n1468) );
    znd3b U497 ( .A(ASKREPLY), .B(n1461), .C(n1595), .Y(n1559) );
    zivb U498 ( .A(n1559), .Y(n1562) );
    zmux21hb U499 ( .A(RXPID[7]), .B(DATA_RX[7]), .S(n1456), .Y(RXPID535_7) );
    zmux21hb U500 ( .A(RXPID[6]), .B(DATA_RX[6]), .S(n1456), .Y(RXPID535_6) );
    zmux21hb U501 ( .A(RXPID[5]), .B(DATA_RX[5]), .S(n1456), .Y(RXPID535_5) );
    zmux21hb U502 ( .A(RXPID[4]), .B(DATA_RX[4]), .S(n1456), .Y(RXPID535_4) );
    zmux21hb U503 ( .A(RXPID[3]), .B(DATA_RX[3]), .S(n1456), .Y(RXPID535_3) );
    zmux21hb U504 ( .A(RXPID[2]), .B(DATA_RX[2]), .S(n1456), .Y(RXPID535_2) );
    zmux21hb U505 ( .A(RXPID[1]), .B(DATA_RX[1]), .S(n1456), .Y(RXPID535_1) );
    zmux21hb U506 ( .A(RXPID[0]), .B(DATA_RX[0]), .S(n1456), .Y(RXPID535_0) );
    zmux21hb U507 ( .A(RXBCNT[10]), .B(RXBCNT981_10), .S(LATCHDAT), .Y(
        RXBCNT989_10) );
    zxo2b U508 ( .A(add_377_carry_10), .B(RXBCNT[10]), .Y(RXBCNT981_10) );
    zmux21hb U509 ( .A(RXBCNT[9]), .B(RXBCNT981_9), .S(LATCHDAT), .Y(
        RXBCNT989_9) );
    zhadrb add_377_U1_1_9 ( .A(RXBCNT[9]), .B(add_377_carry_9), .CO(
        add_377_carry_10), .S(RXBCNT981_9) );
    zmux21hb U510 ( .A(RXBCNT[8]), .B(RXBCNT981_8), .S(LATCHDAT), .Y(
        RXBCNT989_8) );
    zhadrb add_377_U1_1_8 ( .A(RXBCNT[8]), .B(add_377_carry_8), .CO(
        add_377_carry_9), .S(RXBCNT981_8) );
    zmux21hb U511 ( .A(RXBCNT[7]), .B(RXBCNT981_7), .S(LATCHDAT), .Y(
        RXBCNT989_7) );
    zhadrb add_377_U1_1_7 ( .A(RXBCNT[7]), .B(add_377_carry_7), .CO(
        add_377_carry_8), .S(RXBCNT981_7) );
    zmux21hb U512 ( .A(RXBCNT[6]), .B(RXBCNT981_6), .S(LATCHDAT), .Y(
        RXBCNT989_6) );
    zhadrb add_377_U1_1_6 ( .A(RXBCNT[6]), .B(add_377_carry_6), .CO(
        add_377_carry_7), .S(RXBCNT981_6) );
    zmux21hb U513 ( .A(RXBCNT[5]), .B(RXBCNT981_5), .S(LATCHDAT), .Y(
        RXBCNT989_5) );
    zhadrb add_377_U1_1_5 ( .A(RXBCNT[5]), .B(add_377_carry_5), .CO(
        add_377_carry_6), .S(RXBCNT981_5) );
    zmux21hb U514 ( .A(RXBCNT[4]), .B(RXBCNT981_4), .S(LATCHDAT), .Y(
        RXBCNT989_4) );
    zhadrb add_377_U1_1_4 ( .A(RXBCNT[4]), .B(add_377_carry_4), .CO(
        add_377_carry_5), .S(RXBCNT981_4) );
    zmux21hb U515 ( .A(RXBCNT[3]), .B(RXBCNT981_3), .S(LATCHDAT), .Y(
        RXBCNT989_3) );
    zhadrb add_377_U1_1_3 ( .A(RXBCNT[3]), .B(add_377_carry_3), .CO(
        add_377_carry_4), .S(RXBCNT981_3) );
    zmux21hb U516 ( .A(RXBCNT[2]), .B(RXBCNT981_2), .S(LATCHDAT), .Y(
        RXBCNT989_2) );
    zhadrb add_377_U1_1_2 ( .A(RXBCNT[2]), .B(add_377_carry_2), .CO(
        add_377_carry_3), .S(RXBCNT981_2) );
    zmux21hb U517 ( .A(RXBCNT[1]), .B(RXBCNT981_1), .S(LATCHDAT), .Y(
        RXBCNT989_1) );
    zhadrb add_377_U1_1_1 ( .A(RXBCNT[1]), .B(RXBCNT[0]), .CO(add_377_carry_2), 
        .S(RXBCNT981_1) );
    zoai21b U518 ( .A(n1457), .B(n1550), .C(n1551), .Y(ADDSEL1101_0) );
    zmux21hb U519 ( .A(RXADDRF[8]), .B(DATA_RX[0]), .S(n1591), .Y(n_2277) );
    zmux21hb U520 ( .A(RXADDRF[2]), .B(DATA_RX[2]), .S(n1592), .Y(n_1870) );
    zmux21hb U521 ( .A(RXADDRF[12]), .B(DATA_RX[4]), .S(n1591), .Y(n_2269) );
    zmux21hb U522 ( .A(RXADDRF[15]), .B(DATA_RX[7]), .S(n1591), .Y(n_2263) );
    zmux21hb U523 ( .A(RXADDRF[5]), .B(DATA_RX[5]), .S(n1592), .Y(n_1864) );
    zivb U524 ( .A(n1577), .Y(n1569) );
    zivb U525 ( .A(n1563), .Y(n1542) );
    zor2b U526 ( .A(RXACTIVE_SYNC), .B(n1585), .Y(n1563) );
    zivb U527 ( .A(n1545), .Y(n1556) );
    zivb U528 ( .A(EN_CHKTOGCRC), .Y(n1565) );
    zmux21hb U529 ( .A(RXADDRF[21]), .B(DATA_RX[5]), .S(n1590), .Y(n_2670) );
    zmux21hb U530 ( .A(RXADDRF[4]), .B(DATA_RX[4]), .S(n1592), .Y(n_1866) );
    zmux21hb U531 ( .A(RXADDRF[14]), .B(DATA_RX[6]), .S(n1591), .Y(n_2265) );
    zmux21hb U532 ( .A(RXADDRF[20]), .B(DATA_RX[4]), .S(n1590), .Y(n_2672) );
    zdffqrb_ BABBLE_reg ( .CK(CLK60M), .D(BABBLE1031), .R(STSRST_), .Q(BABBLE)
         );
    zmux21hb U533 ( .A(RXADDRF[9]), .B(DATA_RX[1]), .S(n1591), .Y(n_2275) );
    zoai21b U534 ( .A(n1457), .B(n1552), .C(n1553), .Y(ADDSEL1101_1) );
    zmux21hb U535 ( .A(RXADDRF[13]), .B(DATA_RX[5]), .S(n1591), .Y(n_2267) );
    zmux21hb U536 ( .A(RXADDRF[3]), .B(DATA_RX[3]), .S(n1592), .Y(n_1868) );
    zor2b U537 ( .A(n1540), .B(RXACTIVE), .Y(RXACTIVE_SYNC) );
    zan3b U538 ( .A(RVLD_SYNC), .B(RXACTIVE_FLAG), .C(EN_REF_RVLD), .Y(n1540)
         );
    zivb U539 ( .A(RXACTIVE_SYNC), .Y(n1580) );
    zmux21hb U540 ( .A(RXADDRF[19]), .B(DATA_RX[3]), .S(n1590), .Y(n_2674) );
    zmux21hb U541 ( .A(RXADDRF[1]), .B(DATA_RX[1]), .S(n1592), .Y(n_1872) );
    zmux21hb U542 ( .A(RXADDRF[11]), .B(DATA_RX[3]), .S(n1591), .Y(n_2271) );
    zaoi21b U543 ( .A(n1584), .B(n1470), .C(n1461), .Y(CRCEN_T624) );
    zivb U544 ( .A(n1544), .Y(n1470) );
    znd2b U545 ( .A(n1462), .B(n1463), .Y(n1544) );
    zmux21hb U546 ( .A(RXADDRF[17]), .B(DATA_RX[1]), .S(n1590), .Y(n_2678) );
    zmux21hb U547 ( .A(RXADDRF[6]), .B(DATA_RX[6]), .S(n1592), .Y(n_1862) );
    zmux21hb U548 ( .A(RXADDRF[22]), .B(DATA_RX[6]), .S(n1590), .Y(n_2668) );
    zmux21hb U549 ( .A(RXADDRF[7]), .B(DATA_RX[7]), .S(n1592), .Y(n_1860) );
    znr2b U550 ( .A(n1536), .B(n1471), .Y(LATCHDAT783) );
    znd2b U551 ( .A(EN_LATCHDAT), .B(LATCHDAT_P), .Y(n1471) );
    zmux21hb U552 ( .A(RXADDRF[16]), .B(DATA_RX[0]), .S(n1590), .Y(n_2680) );
    zmux21hb U553 ( .A(RXADDRF[23]), .B(DATA_RX[7]), .S(n1590), .Y(n_2666) );
    zmux21hb U554 ( .A(RXADDRF[18]), .B(DATA_RX[2]), .S(n1590), .Y(n_2676) );
    zivb U555 ( .A(n1551), .Y(n1590) );
    znd2b U556 ( .A(n1539), .B(n1457), .Y(n1551) );
    zao21b U557 ( .A(n1541), .B(ASKREPLY), .C(PHYERR), .Y(PHYERR291) );
    zoai21b U558 ( .A(n1457), .B(n1554), .C(n1555), .Y(ADDSEL1101_2) );
    zmux21hb U559 ( .A(RXADDRF[10]), .B(DATA_RX[2]), .S(n1591), .Y(n_2273) );
    zivb U560 ( .A(n1555), .Y(n1591) );
    znd2b U561 ( .A(n1538), .B(n1457), .Y(n1555) );
    zmux21hb U562 ( .A(RXADDRF[0]), .B(DATA_RX[0]), .S(n1592), .Y(n_1874) );
    zivb U563 ( .A(n1553), .Y(n1592) );
    znd2b U564 ( .A(n1537), .B(n1457), .Y(n1553) );
    zan2b U565 ( .A(n1548), .B(RXSM_4), .Y(LATCHADDR) );
    zivb U566 ( .A(n1543), .Y(n1548) );
    zao33b U567 ( .A(RXSM_4), .B(n1558), .C(n1452), .D(RXTOKEN), .E(n1581), 
        .F(n1453), .Y(n1543) );
    zivb U568 ( .A(RXSOF), .Y(n1581) );
    znr2b U569 ( .A(n1536), .B(n1465), .Y(SPD) );
    znd2b U570 ( .A(n1531), .B(n1530), .Y(n1465) );
    zivb U571 ( .A(n1571), .Y(TOGMATCH) );
    zivb U572 ( .A(n1582), .Y(NORMPKT) );
    zcxi7b U573 ( .A(n1546), .B(RXSM_2), .C(RXTOKENPHASE), .D(PKRVEND_T), .E(
        n1547), .Y(PKRVEND) );
    zoai21b U574 ( .A(TMOUT), .B(EOF2), .C(n1594), .Y(n1546) );
    zivb U575 ( .A(RXVALID_SYNC_T), .Y(n1534) );
    zdffqrb RXSM_reg_4 ( .CK(CLK60M), .D(RXSM457_4), .R(TRST_), .Q(RXSM_4) );
    zivb U576 ( .A(RXSM_4), .Y(n1549) );
    zdffqrb RXSM_reg_3 ( .CK(CLK60M), .D(RXSM457_3), .R(TRST_), .Q(RXSM_3) );
    zivb U577 ( .A(RXSM_3), .Y(n1564) );
    zdffqrb RXSM_reg_2 ( .CK(CLK60M), .D(RXSM457_2), .R(TRST_), .Q(RXSM_2) );
    zivb U578 ( .A(RXSM_2), .Y(n1584) );
    zdffqrb RXSM_reg_1 ( .CK(CLK60M), .D(RXSM457_1), .R(TRST_), .Q(RXSM_1) );
    zivb U579 ( .A(RXSM_1), .Y(n1560) );
    zdffqrb RXSM_reg_0 ( .CK(CLK60M), .D(RXSM457_0), .R(TRST_), .Q(RXSM_0) );
    zivb U580 ( .A(RXSM_0), .Y(n1558) );
    zdffqrb HOLD_reg_23 ( .CK(CLK60M), .D(DATA_RX[7]), .R(TRST_), .Q(RXCRCDAT
        [7]) );
    zdffqrb HOLD_reg_22 ( .CK(CLK60M), .D(DATA_RX[6]), .R(TRST_), .Q(RXCRCDAT
        [6]) );
    zdffqrb HOLD_reg_21 ( .CK(CLK60M), .D(DATA_RX[5]), .R(TRST_), .Q(RXCRCDAT
        [5]) );
    zdffqrb HOLD_reg_20 ( .CK(CLK60M), .D(DATA_RX[4]), .R(TRST_), .Q(RXCRCDAT
        [4]) );
    zdffqrb HOLD_reg_19 ( .CK(CLK60M), .D(DATA_RX[3]), .R(TRST_), .Q(RXCRCDAT
        [3]) );
    zdffqrb HOLD_reg_18 ( .CK(CLK60M), .D(DATA_RX[2]), .R(TRST_), .Q(RXCRCDAT
        [2]) );
    zdffqrb HOLD_reg_17 ( .CK(CLK60M), .D(DATA_RX[1]), .R(TRST_), .Q(RXCRCDAT
        [1]) );
    zdffqrb HOLD_reg_16 ( .CK(CLK60M), .D(DATA_RX[0]), .R(TRST_), .Q(RXCRCDAT
        [0]) );
    zdffqrb HOLD_reg_15 ( .CK(CLK60M), .D(n1622), .R(TRST_), .Q(HOLD_15) );
    zdffqrb HOLD_reg_14 ( .CK(CLK60M), .D(n1621), .R(TRST_), .Q(HOLD_14) );
    zdffqrb HOLD_reg_13 ( .CK(CLK60M), .D(n1620), .R(TRST_), .Q(HOLD_13) );
    zdffqrb HOLD_reg_12 ( .CK(CLK60M), .D(n1619), .R(TRST_), .Q(HOLD_12) );
    zdffqrb HOLD_reg_11 ( .CK(CLK60M), .D(n1618), .R(TRST_), .Q(HOLD_11) );
    zdffqrb HOLD_reg_10 ( .CK(CLK60M), .D(n1617), .R(TRST_), .Q(HOLD_10) );
    zdffqrb HOLD_reg_9 ( .CK(CLK60M), .D(n1616), .R(TRST_), .Q(HOLD_9) );
    zdffqrb HOLD_reg_8 ( .CK(CLK60M), .D(n1615), .R(TRST_), .Q(HOLD_8) );
    zdffqrb HOLD_reg_7 ( .CK(CLK60M), .D(n1614), .R(TRST_), .Q(USBDAT[7]) );
    zdffqrb HOLD_reg_6 ( .CK(CLK60M), .D(n1612), .R(TRST_), .Q(USBDAT[6]) );
    zdffqrb HOLD_reg_5 ( .CK(CLK60M), .D(n1610), .R(TRST_), .Q(USBDAT[5]) );
    zdffqrb HOLD_reg_4 ( .CK(CLK60M), .D(n1608), .R(TRST_), .Q(USBDAT[4]) );
    zdffqrb HOLD_reg_3 ( .CK(CLK60M), .D(n1606), .R(TRST_), .Q(USBDAT[3]) );
    zdffqrb HOLD_reg_2 ( .CK(CLK60M), .D(n1604), .R(TRST_), .Q(USBDAT[2]) );
    zdffqrb HOLD_reg_1 ( .CK(CLK60M), .D(n1602), .R(TRST_), .Q(USBDAT[1]) );
    zdffqrb HOLD_reg_0 ( .CK(CLK60M), .D(n1600), .R(TRST_), .Q(USBDAT[0]) );
    zdffqrb RXPID_reg_7 ( .CK(CLK60M), .D(RXPID535_7), .R(STSRST_), .Q(RXPID
        [7]) );
    zdffqrb RXPID_reg_6 ( .CK(CLK60M), .D(RXPID535_6), .R(STSRST_), .Q(RXPID
        [6]) );
    zdffqrb RXPID_reg_5 ( .CK(CLK60M), .D(RXPID535_5), .R(STSRST_), .Q(RXPID
        [5]) );
    zdffqrb RXPID_reg_4 ( .CK(CLK60M), .D(RXPID535_4), .R(STSRST_), .Q(RXPID
        [4]) );
    zdffqrb RXPID_reg_3 ( .CK(CLK60M), .D(RXPID535_3), .R(STSRST_), .Q(RXPID
        [3]) );
    zdffqrb RXPID_reg_2 ( .CK(CLK60M), .D(RXPID535_2), .R(STSRST_), .Q(RXPID
        [2]) );
    zdffqrb RXPID_reg_1 ( .CK(CLK60M), .D(RXPID535_1), .R(STSRST_), .Q(RXPID
        [1]) );
    zdffqrb RXPID_reg_0 ( .CK(CLK60M), .D(RXPID535_0), .R(STSRST_), .Q(RXPID
        [0]) );
    zdffqrb RXBCNT_reg_10 ( .CK(CLK60M), .D(RXBCNT989_10), .R(STSRST_), .Q(
        RXBCNT[10]) );
    zivb U581 ( .A(RXBCNT[10]), .Y(n1483) );
    zdffqrb RXBCNT_reg_9 ( .CK(CLK60M), .D(RXBCNT989_9), .R(STSRST_), .Q(
        RXBCNT[9]) );
    zivb U582 ( .A(RXBCNT[9]), .Y(n1481) );
    zdffqrb RXBCNT_reg_8 ( .CK(CLK60M), .D(RXBCNT989_8), .R(STSRST_), .Q(
        RXBCNT[8]) );
    zivb U583 ( .A(RXBCNT[8]), .Y(n1475) );
    zdffqrb RXBCNT_reg_7 ( .CK(CLK60M), .D(RXBCNT989_7), .R(STSRST_), .Q(
        RXBCNT[7]) );
    zivb U584 ( .A(RXBCNT[7]), .Y(n1473) );
    zdffqrb RXBCNT_reg_6 ( .CK(CLK60M), .D(RXBCNT989_6), .R(STSRST_), .Q(
        RXBCNT[6]) );
    zivb U585 ( .A(RXBCNT[6]), .Y(n1474) );
    zdffqrb RXBCNT_reg_5 ( .CK(CLK60M), .D(RXBCNT989_5), .R(STSRST_), .Q(
        RXBCNT[5]) );
    zivb U586 ( .A(RXBCNT[5]), .Y(n1479) );
    zdffqrb RXBCNT_reg_4 ( .CK(CLK60M), .D(RXBCNT989_4), .R(STSRST_), .Q(
        RXBCNT[4]) );
    zivb U587 ( .A(RXBCNT[4]), .Y(n1477) );
    zdffqrb RXBCNT_reg_3 ( .CK(CLK60M), .D(RXBCNT989_3), .R(STSRST_), .Q(
        RXBCNT[3]) );
    zivb U588 ( .A(RXBCNT[3]), .Y(n1480) );
    zdffqrb RXBCNT_reg_2 ( .CK(CLK60M), .D(RXBCNT989_2), .R(STSRST_), .Q(
        RXBCNT[2]) );
    zivb U589 ( .A(RXBCNT[2]), .Y(n1478) );
    zdffqrb RXBCNT_reg_1 ( .CK(CLK60M), .D(RXBCNT989_1), .R(STSRST_), .Q(
        RXBCNT[1]) );
    zivb U590 ( .A(RXBCNT[1]), .Y(n1476) );
    zdffsb ADDSEL_reg_0 ( .CK(CLK60M), .D(ADDSEL1101_0), .S(STSRST_), .Q(n1537
        ), .QN(n1550) );
    zdffqrb RXADDRF_reg2_8 ( .CK(CLK60M), .D(n_2277), .R(STSRST_), .Q(RXADDRF
        [8]) );
    zdffqrb_ RXCRCRST_reg ( .CK(CLK60M), .D(RXSM_1), .R(TRST_), .Q(RXCRCRST)
         );
    zdffqrb RXADDRF_reg_2 ( .CK(CLK60M), .D(n_1870), .R(STSRST_), .Q(RXADDRF
        [2]) );
    zdffqrb RXADDRF_reg2_12 ( .CK(CLK60M), .D(n_2269), .R(STSRST_), .Q(RXADDRF
        [12]) );
    zdffqrb LATCHPID_reg ( .CK(CLK60M), .D(n1456), .R(STSRST_), .Q(LATCHPID)
         );
    zdffqrb RXVALID_L2H_reg ( .CK(CLK60M), .D(n1598), .R(STSRST_), .Q(
        RXVALID_L2H) );
    zivb U591 ( .A(RXVALID_L2H), .Y(n1467) );
    zdffqrb_ CRCHK_reg ( .CK(CLK60M), .D(RXSM_3), .R(STSRST_), .Q(CRCHK) );
    zdffqrb PKRVEND_T_reg ( .CK(CLK60M), .D(n1597), .R(TRST_), .Q(PKRVEND_T)
         );
    zdffqrb RXADDRF_reg2_15 ( .CK(CLK60M), .D(n_2263), .R(STSRST_), .Q(RXADDRF
        [15]) );
    zdffqrb RXADDRF_reg_5 ( .CK(CLK60M), .D(n_1864), .R(STSRST_), .Q(RXADDRF
        [5]) );
    zdffqrb RXSTART_reg ( .CK(CLK60M), .D(RXSTART587), .R(TRST_), .Q(RXSTART)
         );
    zivb U592 ( .A(RXSTART), .Y(n1547) );
    zdffqrb_ LATCHDAT_P_reg ( .CK(CLK60M), .D(n1596), .R(TRST_), .Q(LATCHDAT_P
        ) );
    zivb U593 ( .A(LATCHDAT_P), .Y(n1494) );
    zdffqrb_ RXCRCEN_reg ( .CK(CLK60M), .D(CRCEN_T), .R(TRST_), .Q(RXCRCEN) );
    zdffqrb RXADDRF_reg3_21 ( .CK(CLK60M), .D(n_2670), .R(STSRST_), .Q(RXADDRF
        [21]) );
    zdffqrb RXADDRF_reg_4 ( .CK(CLK60M), .D(n_1866), .R(STSRST_), .Q(RXADDRF
        [4]) );
    zdffqrb RXADDRF_reg2_14 ( .CK(CLK60M), .D(n_2265), .R(STSRST_), .Q(RXADDRF
        [14]) );
    zdffqrb RXADDRF_reg3_20 ( .CK(CLK60M), .D(n_2672), .R(STSRST_), .Q(RXADDRF
        [20]) );
    zdffqrb RXADDRF_reg2_9 ( .CK(CLK60M), .D(n_2275), .R(STSRST_), .Q(RXADDRF
        [9]) );
    zdffrb ADDSEL_reg_1 ( .CK(CLK60M), .D(ADDSEL1101_1), .R(STSRST_), .Q(n1538
        ), .QN(n1552) );
    zdffqrb RXADDRF_reg2_13 ( .CK(CLK60M), .D(n_2267), .R(STSRST_), .Q(RXADDRF
        [13]) );
    zdffqrb RXADDRF_reg_3 ( .CK(CLK60M), .D(n_1868), .R(STSRST_), .Q(RXADDRF
        [3]) );
    zdffqrb RXACTIVE_FLAG_reg ( .CK(CLK60M), .D(RXACTIVE_SYNC), .R(STSRST_), 
        .Q(RXACTIVE_FLAG) );
    zdffqrb RXADDRF_reg3_19 ( .CK(CLK60M), .D(n_2674), .R(STSRST_), .Q(RXADDRF
        [19]) );
    zdffqrb RXADDRF_reg_1 ( .CK(CLK60M), .D(n_1872), .R(STSRST_), .Q(RXADDRF
        [1]) );
    zdffqrb RXADDRF_reg2_11 ( .CK(CLK60M), .D(n_2271), .R(STSRST_), .Q(RXADDRF
        [11]) );
    zdffqrb CRCEN_T_reg ( .CK(CLK60M), .D(CRCEN_T624), .R(TRST_), .Q(CRCEN_T)
         );
    zdffqrb RXADDRF_reg3_17 ( .CK(CLK60M), .D(n_2678), .R(STSRST_), .Q(RXADDRF
        [17]) );
    zdffqrb RVLD_SYNC_reg ( .CK(CLK60M), .D(RVLD), .R(STSRST_), .Q(RVLD_SYNC)
         );
    zdffqrb_ RXVALID_SYNC_2T_reg ( .CK(CLK60M), .D(RXVALID), .R(STSRST_), .Q(
        RXVALID_SYNC_2T) );
    zivb U594 ( .A(RXVALID_SYNC_2T), .Y(n1535) );
    zdffqrb RXADDRF_reg_6 ( .CK(CLK60M), .D(n_1862), .R(STSRST_), .Q(RXADDRF
        [6]) );
    zdffqrb RXADDRF_reg3_22 ( .CK(CLK60M), .D(n_2668), .R(STSRST_), .Q(RXADDRF
        [22]) );
    zdffqrb RXADDRF_reg_7 ( .CK(CLK60M), .D(n_1860), .R(STSRST_), .Q(RXADDRF
        [7]) );
    zdffqrb_ LATCHDAT_reg ( .CK(CLK60M), .D(LATCHDAT783), .R(TRST_), .Q(
        LATCHDAT) );
    zdffqrb RXADDRF_reg3_16 ( .CK(CLK60M), .D(n_2680), .R(STSRST_), .Q(RXADDRF
        [16]) );
    zdffqrb RXADDRF_reg3_23 ( .CK(CLK60M), .D(n_2666), .R(STSRST_), .Q(RXADDRF
        [23]) );
    zdffqrb RXADDRF_reg3_18 ( .CK(CLK60M), .D(n_2676), .R(STSRST_), .Q(RXADDRF
        [18]) );
    zdffqrb PHYERR_reg ( .CK(CLK60M), .D(PHYERR291), .R(STSRST_), .Q(PHYERR)
         );
    zivb U595 ( .A(PHYERR), .Y(n1574) );
    zdffrb ADDSEL_reg_2 ( .CK(CLK60M), .D(ADDSEL1101_2), .R(STSRST_), .Q(n1539
        ), .QN(n1554) );
    zdffqrb RXADDRF_reg2_10 ( .CK(CLK60M), .D(n_2273), .R(STSRST_), .Q(RXADDRF
        [10]) );
    zdffqrb RXADDRF_reg_0 ( .CK(CLK60M), .D(n_1874), .R(STSRST_), .Q(RXADDRF
        [0]) );
    znr5b U596 ( .A(RXSM_1), .B(RXSM_3), .C(RXSM_2), .D(n1580), .E(n1577), .Y(
        n1452) );
    znr4b U597 ( .A(n1576), .B(n1577), .C(PIDERR), .D(n1455), .Y(n1453) );
    znr2b U598 ( .A(RXSM_0), .B(n1574), .Y(n1454) );
    zan3b U599 ( .A(DATAIN), .B(n1565), .C(n1571), .Y(n1455) );
    zivb U600 ( .A(RXBCNT[0]), .Y(RXBCNT981_0) );
    zdffqrb RXBCNT_reg_0 ( .CK(CLK60M), .D(RXBCNT989_0), .R(STSRST_), .Q(
        RXBCNT[0]) );
    zivb U601 ( .A(RXDATA), .Y(n1573) );
    zan3b U602 ( .A(n1493), .B(n1594), .C(n1569), .Y(n1456) );
    znd2b U603 ( .A(ASKREPLY), .B(n1469), .Y(n1557) );
    zivb U604 ( .A(n1557), .Y(n1561) );
    znd2b U605 ( .A(n1560), .B(n1464), .Y(n1583) );
    zivb U606 ( .A(n1583), .Y(n1594) );
    zoa21d U607 ( .A(RXSM_4), .B(n1543), .C(RXVALID), .Y(n1457) );
    ziv11b U608 ( .A(MAXLEN[10]), .Y(n1459), .Z(n1458) );
    zivb U609 ( .A(n1461), .Y(n1460) );
    zivb U610 ( .A(RXVALID), .Y(n1461) );
    zao21d U611 ( .A(n1466), .B(n1467), .C(RXVALID), .Y(EN_LATCHDAT) );
    zivh U614 ( .A(MAXLEN[7]), .Y(n1484) );
    zivh U615 ( .A(MAXLEN[6]), .Y(n1485) );
    zivh U616 ( .A(MAXLEN[8]), .Y(n1486) );
    zivh U617 ( .A(MAXLEN[1]), .Y(n1487) );
    zivh U618 ( .A(MAXLEN[4]), .Y(n1488) );
    zivh U619 ( .A(MAXLEN[5]), .Y(n1490) );
    zivh U620 ( .A(MAXLEN[3]), .Y(n1491) );
    zivh U621 ( .A(MAXLEN[9]), .Y(n1492) );
    znd2d U622 ( .A(n1496), .B(n1497), .Y(n1495) );
    znd2d U623 ( .A(n1499), .B(n1500), .Y(n1498) );
    znd3d U624 ( .A(n1502), .B(RXBCNT981_0), .C(n1503), .Y(n1501) );
    zan6d U625 ( .A(n1504), .B(n1505), .C(n1506), .D(n1507), .E(n1508), .F(
        n1509), .Y(n1500) );
    zan5d U626 ( .A(n1510), .B(n1511), .C(n1512), .D(n1513), .E(n1514), .Y(
        n1499) );
    znr3d U627 ( .A(n1494), .B(MAC_SLAVE_ACT), .C(n1532), .Y(n1472) );
    znd2d U628 ( .A(RXBCNT[10]), .B(n1459), .Y(n1507) );
    znd2d U629 ( .A(MAXLEN[7]), .B(n1473), .Y(n1509) );
    znd2d U630 ( .A(MAXLEN[6]), .B(n1474), .Y(n1505) );
    znd2d U631 ( .A(MAXLEN[8]), .B(n1475), .Y(n1504) );
    znd2d U632 ( .A(MAXLEN[1]), .B(n1476), .Y(n1506) );
    znd2d U633 ( .A(MAXLEN[4]), .B(n1477), .Y(n1511) );
    znd2d U634 ( .A(MAXLEN[5]), .B(n1479), .Y(n1512) );
    znd2d U635 ( .A(MAXLEN[3]), .B(n1480), .Y(n1514) );
    znd2d U636 ( .A(MAXLEN[9]), .B(n1481), .Y(n1513) );
    znd2d U637 ( .A(RXBCNT[6]), .B(n1485), .Y(n1521) );
    znd2d U638 ( .A(RXBCNT[8]), .B(n1486), .Y(n1520) );
    znd2d U639 ( .A(RXBCNT[1]), .B(n1487), .Y(n1522) );
    znd2d U640 ( .A(RXBCNT[4]), .B(n1488), .Y(n1525) );
    znd2d U641 ( .A(RXBCNT[5]), .B(n1490), .Y(n1526) );
    znd2d U642 ( .A(RXBCNT[3]), .B(n1491), .Y(n1529) );
    znd2d U643 ( .A(RXBCNT[9]), .B(n1492), .Y(n1528) );
    zmux21ld U644 ( .A(n1498), .B(n1501), .S(MAC_SLAVE_ACT), .Y(n1497) );
    zivl U645 ( .A(n1495), .Y(n1536) );
    zdffqrb RXVALID_SYNC_T_reg ( .CK(CLK60M), .D(n1460), .R(STSRST_), .Q(
        RXVALID_SYNC_T) );
    zor6b U646 ( .A(RXACTIVE_SYNC), .B(n1456), .C(n1542), .D(n1543), .E(n1544), 
        .F(n1545), .Y(RXSTART587) );
    zoai22d U647 ( .A(n1556), .B(n1557), .C(n1558), .D(n1559), .Y(RXSM457_0)
         );
    zoai22d U648 ( .A(n1557), .B(n1563), .C(n1559), .D(n1564), .Y(RXSM457_3)
         );
    zoai22d U649 ( .A(n1548), .B(n1557), .C(n1549), .D(n1559), .Y(RXSM457_4)
         );
    zmux21ld U651 ( .A(n1572), .B(SL_TOGMATCH), .S(MAC_SLAVE_ACT), .Y(n1571)
         );
    zor3b U652 ( .A(RXSM_3), .B(RXSM_0), .C(RXSM_4), .Y(n1575) );
    zor3b U653 ( .A(RXSM_2), .B(n1560), .C(n1575), .Y(n1576) );
    zor4b U654 ( .A(PHYERR), .B(BABBLE), .C(CRCERR), .D(PIDERR), .Y(n1582) );
    zor3b U655 ( .A(n1584), .B(n1583), .C(n1577), .Y(n1585) );
    zao211b U656 ( .A(n1454), .B(n1586), .C(n1566), .D(n1567), .Y(n1545) );
    zoai21d U657 ( .A(n1573), .B(n1588), .C(n1589), .Y(n1572) );
    zind2d U658 ( .A(EXEITD), .B(ISO), .Y(n1588) );
    zaoi2x4d U659 ( .A(DAT1), .B(RXDATA1), .C(DAT0), .D(RXDATA0), .E(DAT2), 
        .F(RXDATA2), .G(DATM), .H(RXMDATA), .Y(n1589) );
    zor3b U660 ( .A(RXHAND), .B(RXSOF), .C(PIDERR), .Y(n1593) );
    zinr2b U661 ( .A(RXEOPERR), .B(DISCHKEOPERR), .Y(n1541) );
    zao211b U662 ( .A(n1579), .B(n1573), .C(n1593), .D(n1455), .Y(n1570) );
    zbfb U663 ( .A(val832_1), .Y(n1596) );
    zoa21b U664 ( .A(TOGMATCH), .B(n1565), .C(RXCRCEN), .Y(val832_1) );
    zbfb U665 ( .A(RXSTART), .Y(n1597) );
    zbfb U666 ( .A(RXVALID_L2H736), .Y(n1598) );
    zinr2d U667 ( .A(RXVALID), .B(RXVALID_SYNC_T), .Y(RXVALID_L2H736) );
    zivb U668 ( .A(HOLD_8), .Y(n1599) );
    zivb U669 ( .A(n1599), .Y(n1600) );
    zivb U670 ( .A(HOLD_9), .Y(n1601) );
    zivb U671 ( .A(n1601), .Y(n1602) );
    zivb U672 ( .A(HOLD_10), .Y(n1603) );
    zivb U673 ( .A(n1603), .Y(n1604) );
    zivb U674 ( .A(HOLD_11), .Y(n1605) );
    zivb U675 ( .A(n1605), .Y(n1606) );
    zivb U676 ( .A(HOLD_12), .Y(n1607) );
    zivb U677 ( .A(n1607), .Y(n1608) );
    zivb U678 ( .A(HOLD_13), .Y(n1609) );
    zivb U679 ( .A(n1609), .Y(n1610) );
    zivb U680 ( .A(HOLD_14), .Y(n1611) );
    zivb U681 ( .A(n1611), .Y(n1612) );
    zivb U682 ( .A(HOLD_15), .Y(n1613) );
    zivb U683 ( .A(n1613), .Y(n1614) );
    zbfb U684 ( .A(RXCRCDAT[0]), .Y(n1615) );
    zbfb U685 ( .A(RXCRCDAT[1]), .Y(n1616) );
    zbfb U686 ( .A(RXCRCDAT[2]), .Y(n1617) );
    zbfb U687 ( .A(RXCRCDAT[3]), .Y(n1618) );
    zbfb U688 ( .A(RXCRCDAT[4]), .Y(n1619) );
    zbfb U689 ( .A(RXCRCDAT[5]), .Y(n1620) );
    zbfb U690 ( .A(RXCRCDAT[6]), .Y(n1621) );
    zbfb U691 ( .A(RXCRCDAT[7]), .Y(n1622) );
    zao21b U692 ( .A(n1472), .B(n1536), .C(BABBLE), .Y(BABBLE1031) );
endmodule


module HS_CRC ( DATAIN, ADRENDPS, CRC, CRC16, CLK60M, CRCEN, CRCRST, SPLIT, 
    CRCHK, STSRST_, RXDATA, CRCERR, MAC_SLAVE_ACT, SL_CRC16 );
input  [7:0] DATAIN;
input  [18:0] ADRENDPS;
output [15:0] CRC;
input  [15:0] SL_CRC16;
input  CRC16, CLK60M, CRCEN, CRCRST, SPLIT, CRCHK, STSRST_, RXDATA, 
    MAC_SLAVE_ACT;
output CRCERR;
    wire CRCREG_5, C13, PKTCRC16_12, SPAREO6, PKTCRC16298_14, CRCHOLD224_5, 
        PKTCRC16298_7, CRCREG199_15, CRCHOLD224_14, CRCREG199_0, CRCHOLD_16, 
        h7, PKTCRC16_2, CRCREG199_9, PKTCRC16298_9, PKTCRC16_5, h0, CRCHOLD_11, 
        SPAREO0_, CRCREG_2, SPAREO8, CRCREG199_12, C9, PKTCRC16298_0, 
        CRCHOLD224_2, CRCERR128, CRCSFT235_2, CRCREG199_7, CRCHOLD224_13, 
        PKTCRC16298_13, C14, CRCHOLD_18, SPAREO1, PKTCRC16_15, CRCSFT_2, 
        SPAREO9, C15, CRCHOLD_10, h1, PKTCRC16298_8, PKTCRC16_4, PKTCRC16_14, 
        SPAREO0, PKTCRC16298_12, CRCREG_4, CRCREG_3, CRCREG199_13, 
        PKTCRC16298_1, CRCHOLD224_3, n_985, CRCREG199_6, CRCHOLD224_12, 
        CRCHOLD224_4, C12, PKTCRC16298_6, CRCREG199_14, CRCHOLD224_15, 
        CRCREG199_1, PKTCRC16298_15, SPAREO7, PKTCRC16_13, RB11, PKTCRC16_3, 
        CRCREG199_8, CRCHOLD_17, h6, CRCREG_6, C10, SELRC260, PKTCRC16_11, 
        CRCHOLD_8, SPAREO5, PKTCRC16_8, CRCREG199_3, CRCHOLD224_17, 
        CRCHOLD224_6, PKTCRC16298_4, RC13, CRCHOLD_15, CRCREG_8, h4, 
        PKTCRC16_6, RB13, PKTCRC16_1, n_989, RB14, CRCHOLD224_8, h3, 
        CRCHOLD_12, CRCSFT_0, CRCREG_1, RC14, CRCHOLD224_10, CRCREG199_4, 
        n_987, CRCSFT235_1, PKTCRC16298_3, CRCHOLD224_1, CRCREG199_11, 
        PKTCRC16298_10, SPAREO2, RC15, CRCSFT_1, CRCHOLD_13, h2, PKTCRC16_7, 
        RB15, CRCHOLD224_18, CRCHOLD224_9, SPAREO3, SPAREO1_, CRCREG_7, 
        CRCREG_0, PKTCRC16298_11, CRCHOLD224_11, CRCREG199_5, n_986, 
        CRCSFT235_0, PKTCRC16298_2, CRCREG199_10, CRCHOLD224_0, PKTCRC16_9, 
        CRCREG199_2, CRCHOLD224_16, CRCHOLD224_7, C11, PKTCRC16298_5, SPAREO4, 
        CRCHOLD_9, PKTCRC16_10, RB12, n_988, PKTCRC16_0, CRCHOLD_14, h5, n353, 
        n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
        n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
        n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
        n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
        n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
        n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
        n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
        n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
        n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
        n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
        n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
        n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
        n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
        n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
        n553, n554, n555, n556, n557;
    znd3b SPARE629 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE620 ( .CK(CLK60M), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE627 ( .A(SPAREO4), .Y(SPAREO5) );
    znr3b SPARE626 ( .A(SPAREO2), .B(n353), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE628 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE621 ( .CK(1'b0), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zaoi211b SPARE623 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zoai21b SPARE624 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zoai21b SPARE625 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE622 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zmux21hb U144 ( .A(RB11), .B(n389), .S(n353), .Y(n_989) );
    zymx24hb U145 ( .A1(RB15), .A2(RB14), .A3(RB13), .A4(RB12), .B1(RC15), 
        .B2(RC14), .B3(RC13), .B4(n388), .S(n353), .Y1(n_985), .Y2(n_986), 
        .Y3(n_987), .Y4(n_988) );
    zxo2b U146 ( .A(n495), .B(n401), .Y(n494) );
    zxo2b U147 ( .A(n397), .B(n523), .Y(n495) );
    zxo2b U148 ( .A(h4), .B(h5), .Y(n519) );
    zxo2b U149 ( .A(h4), .B(h1), .Y(n521) );
    znd8b U150 ( .A(n535), .B(n536), .C(n537), .D(n538), .E(n539), .F(n540), 
        .G(n541), .H(n542), .Y(n534) );
    zxo2b U151 ( .A(n467), .B(SL_CRC16[7]), .Y(n535) );
    zxo2b U152 ( .A(n468), .B(SL_CRC16[6]), .Y(n536) );
    zxo2b U153 ( .A(n469), .B(SL_CRC16[5]), .Y(n537) );
    zxo2b U154 ( .A(n470), .B(SL_CRC16[4]), .Y(n538) );
    zxo2b U155 ( .A(n471), .B(SL_CRC16[3]), .Y(n539) );
    zxo2b U156 ( .A(n472), .B(SL_CRC16[2]), .Y(n540) );
    zxo2b U157 ( .A(n476), .B(SL_CRC16[1]), .Y(n541) );
    zxo2b U158 ( .A(n477), .B(SL_CRC16[0]), .Y(n542) );
    zxo2b U159 ( .A(PKTCRC16_10), .B(SL_CRC16[10]), .Y(n506) );
    zxo2b U160 ( .A(PKTCRC16_11), .B(SL_CRC16[11]), .Y(n507) );
    zxo2b U161 ( .A(PKTCRC16_8), .B(SL_CRC16[8]), .Y(n504) );
    zxo2b U162 ( .A(PKTCRC16_9), .B(SL_CRC16[9]), .Y(n505) );
    zxo2b U163 ( .A(PKTCRC16_13), .B(SL_CRC16[13]), .Y(n509) );
    zxo2b U164 ( .A(PKTCRC16_12), .B(SL_CRC16[12]), .Y(n508) );
    zxo2b U165 ( .A(PKTCRC16_15), .B(SL_CRC16[15]), .Y(n511) );
    zxo2b U166 ( .A(PKTCRC16_14), .B(SL_CRC16[14]), .Y(n510) );
    zxo2b U167 ( .A(n497), .B(n498), .Y(n496) );
    zxo2b U168 ( .A(n398), .B(n400), .Y(n497) );
    zxo2b U169 ( .A(n525), .B(n494), .Y(n498) );
    zxo2b U170 ( .A(n483), .B(n484), .Y(RB14) );
    zxo2b U171 ( .A(h4), .B(n387), .Y(n483) );
    zxo2b U172 ( .A(n390), .B(n391), .Y(n484) );
    zxo2b U173 ( .A(n485), .B(n486), .Y(RB13) );
    zxo2b U174 ( .A(n392), .B(n519), .Y(n485) );
    zxo2b U175 ( .A(n393), .B(n394), .Y(n486) );
    zivb U176 ( .A(CRC16), .Y(n481) );
    zxo2b U177 ( .A(n488), .B(n489), .Y(RB11) );
    zxo2b U178 ( .A(h2), .B(n521), .Y(n488) );
    zxo2b U179 ( .A(n394), .B(n395), .Y(n489) );
    zxo2b U180 ( .A(DATAIN[3]), .B(DATAIN[4]), .Y(n492) );
    zivb U181 ( .A(DATAIN[4]), .Y(n474) );
    zivb U182 ( .A(DATAIN[7]), .Y(n473) );
    zxo2b U183 ( .A(n528), .B(n529), .Y(n500) );
    zxo2b U184 ( .A(n398), .B(n399), .Y(n528) );
    zxo2b U185 ( .A(n400), .B(n401), .Y(n529) );
    zxo2b U186 ( .A(n397), .B(n527), .Y(n499) );
    zivb U187 ( .A(DATAIN[0]), .Y(n466) );
    zxo2b U188 ( .A(n393), .B(n526), .Y(n527) );
    zxo2b U189 ( .A(n533), .B(n501), .Y(n503) );
    zxo2b U190 ( .A(n531), .B(n532), .Y(n533) );
    zxo2b U191 ( .A(n402), .B(n401), .Y(n501) );
    zxo2b U192 ( .A(CRCREG_1), .B(n396), .Y(n433) );
    zxo2b U193 ( .A(n397), .B(n490), .Y(n431) );
    zxo2b U194 ( .A(n465), .B(n491), .Y(n429) );
    zivb U195 ( .A(DATAIN[1]), .Y(n465) );
    zxo2b U196 ( .A(n398), .B(n399), .Y(n427) );
    zxo2b U197 ( .A(n391), .B(n492), .Y(n425) );
    zxo2b U198 ( .A(n400), .B(n401), .Y(n423) );
    zivf U199 ( .A(n410), .Y(n412) );
    zxo2b U200 ( .A(DATAIN[6]), .B(n493), .Y(n421) );
    zxo2b U201 ( .A(n402), .B(n403), .Y(n419) );
    zxo2b U202 ( .A(n499), .B(n500), .Y(n417) );
    zxo2b U203 ( .A(n502), .B(n503), .Y(n415) );
    zan2b U204 ( .A(n414), .B(n404), .Y(SELRC260) );
    zmux21lb U205 ( .A(n479), .B(n478), .S(SPLIT), .Y(n414) );
    zmux21hb U206 ( .A(CRCERR), .B(n517), .S(CRCHK), .Y(CRCERR128) );
    zmux21hb U207 ( .A(n512), .B(n513), .S(RXDATA), .Y(n517) );
    zdffsb CRCREG_reg_8 ( .CK(CLK60M), .D(CRCREG199_8), .S(STSRST_), .Q(
        CRCREG_8), .QN(CRC[7]) );
    zdffsb CRCREG_reg_7 ( .CK(CLK60M), .D(CRCREG199_7), .S(STSRST_), .Q(
        CRCREG_7), .QN(CRC[8]) );
    zdffsb CRCREG_reg_6 ( .CK(CLK60M), .D(CRCREG199_6), .S(STSRST_), .Q(
        CRCREG_6), .QN(CRC[9]) );
    zdffsb CRCREG_reg_5 ( .CK(CLK60M), .D(CRCREG199_5), .S(STSRST_), .Q(
        CRCREG_5), .QN(CRC[10]) );
    zdffsb CRCREG_reg_4 ( .CK(CLK60M), .D(CRCREG199_4), .S(STSRST_), .Q(
        CRCREG_4), .QN(CRC[11]) );
    zdffsb CRCREG_reg_3 ( .CK(CLK60M), .D(CRCREG199_3), .S(STSRST_), .Q(
        CRCREG_3), .QN(CRC[12]) );
    zdffsb CRCREG_reg_2 ( .CK(CLK60M), .D(CRCREG199_2), .S(STSRST_), .Q(
        CRCREG_2), .QN(CRC[13]) );
    zdffsb CRCREG_reg_1 ( .CK(CLK60M), .D(CRCREG199_1), .S(STSRST_), .Q(
        CRCREG_1), .QN(CRC[14]) );
    zdffsb CRCREG_reg_0 ( .CK(CLK60M), .D(CRCREG199_0), .S(STSRST_), .Q(
        CRCREG_0), .QN(CRC[15]) );
    zdffqb CRCHOLD_reg_18 ( .CK(CLK60M), .D(n557), .Q(CRCHOLD_18) );
    zdffqb CRCHOLD_reg_17 ( .CK(CLK60M), .D(n556), .Q(CRCHOLD_17) );
    zdffqb CRCHOLD_reg_16 ( .CK(CLK60M), .D(n555), .Q(CRCHOLD_16) );
    zdffqb CRCHOLD_reg_15 ( .CK(CLK60M), .D(n554), .Q(CRCHOLD_15) );
    zdffqb CRCHOLD_reg_14 ( .CK(CLK60M), .D(n553), .Q(CRCHOLD_14) );
    zdffqb CRCHOLD_reg_13 ( .CK(CLK60M), .D(n552), .Q(CRCHOLD_13) );
    zdffqb CRCHOLD_reg_12 ( .CK(CLK60M), .D(n551), .Q(CRCHOLD_12) );
    zdffqb CRCHOLD_reg_11 ( .CK(CLK60M), .D(n550), .Q(CRCHOLD_11) );
    zdffqb CRCHOLD_reg_10 ( .CK(CLK60M), .D(CRCHOLD224_10), .Q(CRCHOLD_10) );
    zdffqb CRCHOLD_reg_9 ( .CK(CLK60M), .D(CRCHOLD224_9), .Q(CRCHOLD_9) );
    zdffqb CRCHOLD_reg_8 ( .CK(CLK60M), .D(CRCHOLD224_8), .Q(CRCHOLD_8) );
    zdffqb CRCHOLD_reg_7 ( .CK(CLK60M), .D(CRCHOLD224_7), .Q(h7) );
    zivb U208 ( .A(h7), .Y(n462) );
    zdffqb CRCHOLD_reg_6 ( .CK(CLK60M), .D(CRCHOLD224_6), .Q(h6) );
    zivb U209 ( .A(h6), .Y(n461) );
    zdffqb CRCHOLD_reg_5 ( .CK(CLK60M), .D(CRCHOLD224_5), .Q(h5) );
    zdffqb CRCHOLD_reg_4 ( .CK(CLK60M), .D(CRCHOLD224_4), .Q(h4) );
    zdffqb CRCHOLD_reg_3 ( .CK(CLK60M), .D(CRCHOLD224_3), .Q(h3) );
    zdffqb CRCHOLD_reg_2 ( .CK(CLK60M), .D(CRCHOLD224_2), .Q(h2) );
    zivb U210 ( .A(h2), .Y(n460) );
    zdffqb CRCHOLD_reg_1 ( .CK(CLK60M), .D(CRCHOLD224_1), .Q(h1) );
    zivb U211 ( .A(h1), .Y(n459) );
    zdffqb CRCHOLD_reg_0 ( .CK(CLK60M), .D(CRCHOLD224_0), .Q(h0) );
    zivb U212 ( .A(h0), .Y(n458) );
    zdffqb CRCSFT_reg_2 ( .CK(CLK60M), .D(CRCSFT235_2), .Q(CRCSFT_2) );
    zivb U213 ( .A(CRCSFT_2), .Y(n478) );
    zdffqb CRCSFT_reg_1 ( .CK(CLK60M), .D(CRCSFT235_1), .Q(CRCSFT_1) );
    zivb U214 ( .A(CRCSFT_1), .Y(n479) );
    zdffqb CRCSFT_reg_0 ( .CK(CLK60M), .D(CRCSFT235_0), .Q(CRCSFT_0) );
    zivb U215 ( .A(CRCSFT_0), .Y(n480) );
    zdffqsb PKTCRC16_reg_14 ( .CK(CLK60M), .D(PKTCRC16298_14), .S(STSRST_), 
        .Q(PKTCRC16_14) );
    zdffqsb PKTCRC16_reg_13 ( .CK(CLK60M), .D(PKTCRC16298_13), .S(STSRST_), 
        .Q(PKTCRC16_13) );
    zdffqsb PKTCRC16_reg_12 ( .CK(CLK60M), .D(PKTCRC16298_12), .S(STSRST_), 
        .Q(PKTCRC16_12) );
    zdffqsb PKTCRC16_reg_11 ( .CK(CLK60M), .D(PKTCRC16298_11), .S(STSRST_), 
        .Q(PKTCRC16_11) );
    zdffqsb PKTCRC16_reg_10 ( .CK(CLK60M), .D(PKTCRC16298_10), .S(STSRST_), 
        .Q(PKTCRC16_10) );
    zdffqsb PKTCRC16_reg_8 ( .CK(CLK60M), .D(PKTCRC16298_8), .S(STSRST_), .Q(
        PKTCRC16_8) );
    zdffqsb PKTCRC16_reg_7 ( .CK(CLK60M), .D(PKTCRC16298_7), .S(STSRST_), .Q(
        PKTCRC16_7) );
    zivb U216 ( .A(PKTCRC16_7), .Y(n467) );
    zivb U217 ( .A(PKTCRC16_6), .Y(n468) );
    zivb U218 ( .A(PKTCRC16_5), .Y(n469) );
    zdffqsb PKTCRC16_reg_4 ( .CK(CLK60M), .D(PKTCRC16298_4), .S(STSRST_), .Q(
        PKTCRC16_4) );
    zivb U219 ( .A(PKTCRC16_4), .Y(n470) );
    zivb U220 ( .A(PKTCRC16_3), .Y(n471) );
    zdffqsb PKTCRC16_reg_2 ( .CK(CLK60M), .D(PKTCRC16298_2), .S(STSRST_), .Q(
        PKTCRC16_2) );
    zivb U221 ( .A(PKTCRC16_2), .Y(n472) );
    zdffqsb PKTCRC16_reg_1 ( .CK(CLK60M), .D(PKTCRC16298_1), .S(STSRST_), .Q(
        PKTCRC16_1) );
    zivb U222 ( .A(PKTCRC16_1), .Y(n476) );
    zdffqsb PKTCRC16_reg_0 ( .CK(CLK60M), .D(PKTCRC16298_0), .S(STSRST_), .Q(
        PKTCRC16_0) );
    zivb U223 ( .A(PKTCRC16_0), .Y(n477) );
    zdffqrb_ SELRC_reg ( .CK(CLK60M), .D(SELRC260), .R(STSRST_), .Q(n353) );
    zdffqrb CRCERR_reg ( .CK(CLK60M), .D(CRCERR128), .R(STSRST_), .Q(CRCERR)
         );
    znr2d U224 ( .A(n464), .B(n481), .Y(n385) );
    znr2b U225 ( .A(CRC16), .B(n464), .Y(n386) );
    zxn2b U226 ( .A(n458), .B(C15), .Y(n387) );
    zxn2b U227 ( .A(n459), .B(C14), .Y(n388) );
    zxn2b U228 ( .A(n460), .B(C13), .Y(n389) );
    zxn2b U229 ( .A(n461), .B(h3), .Y(n390) );
    zxn2b U230 ( .A(CRC[3]), .B(C11), .Y(n391) );
    zxn2b U231 ( .A(n459), .B(h0), .Y(n392) );
    zxn2b U232 ( .A(CRC[1]), .B(C15), .Y(n393) );
    zxn2b U233 ( .A(n462), .B(C11), .Y(n394) );
    zxn2b U234 ( .A(CRC[1]), .B(C13), .Y(n395) );
    zxn2b U235 ( .A(n466), .B(C15), .Y(n396) );
    zxn2b U236 ( .A(n466), .B(DATAIN[1]), .Y(n397) );
    zxn2b U237 ( .A(CRC[3]), .B(C13), .Y(n398) );
    zxn2b U238 ( .A(n475), .B(DATAIN[3]), .Y(n399) );
    zxn2b U239 ( .A(CRC[4]), .B(C10), .Y(n400) );
    zxn2b U240 ( .A(n474), .B(DATAIN[5]), .Y(n401) );
    zxn2b U241 ( .A(n473), .B(DATAIN[6]), .Y(n402) );
    zxn2b U242 ( .A(CRC[7]), .B(C9), .Y(n403) );
    ziv11b U243 ( .A(CRCRST), .Y(n404), .Z(n405) );
    zao22b U244 ( .A(CRCHOLD_14), .B(n548), .C(ADRENDPS[14]), .D(n409), .Y(
        CRCHOLD224_14) );
    zao22b U245 ( .A(CRCHOLD_17), .B(n548), .C(ADRENDPS[17]), .D(n405), .Y(
        CRCHOLD224_17) );
    zao22b U246 ( .A(CRCHOLD_11), .B(n548), .C(ADRENDPS[11]), .D(n405), .Y(
        CRCHOLD224_11) );
    zan2b U247 ( .A(n548), .B(CRCREG_2), .Y(n420) );
    zan2b U248 ( .A(n548), .B(CRCREG_5), .Y(n426) );
    zan2b U249 ( .A(n548), .B(CRCREG_8), .Y(n432) );
    ziv22d U250 ( .A(n463), .Y1(n407), .Y2(n406) );
    zivh U251 ( .A(n406), .Y(n408) );
    zao22b U252 ( .A(CRCHOLD_12), .B(n407), .C(ADRENDPS[12]), .D(n409), .Y(
        CRCHOLD224_12) );
    zao22b U253 ( .A(CRCHOLD_15), .B(n408), .C(ADRENDPS[15]), .D(CRCRST), .Y(
        CRCHOLD224_15) );
    zao22b U254 ( .A(CRCHOLD_18), .B(n407), .C(ADRENDPS[18]), .D(n405), .Y(
        CRCHOLD224_18) );
    zan2b U255 ( .A(n407), .B(CRCREG_1), .Y(n418) );
    zan2b U256 ( .A(n549), .B(CRCREG_4), .Y(n424) );
    zan2b U257 ( .A(n549), .B(CRCREG_7), .Y(n430) );
    zivb U258 ( .A(n404), .Y(n409) );
    ziv22d U259 ( .A(n464), .Y1(n411), .Y2(n410) );
    zao22b U260 ( .A(CRCSFT_1), .B(n412), .C(CRCSFT_2), .D(n407), .Y(
        CRCSFT235_2) );
    zan2b U261 ( .A(n412), .B(PKTCRC16_9), .Y(n443) );
    znd2d U262 ( .A(n404), .B(n413), .Y(n464) );
    ziv13d U263 ( .A(CRCEN), .Y2(n413) );
    zivb U264 ( .A(n404), .Y(n546) );
    zdffsd CRCREG_reg_15 ( .CK(CLK60M), .D(CRCREG199_15), .S(STSRST_), .Q(C15), 
        .QN(CRC[0]) );
    zdffsd CRCREG_reg_14 ( .CK(CLK60M), .D(CRCREG199_14), .S(STSRST_), .Q(C14), 
        .QN(CRC[1]) );
    zdffsd CRCREG_reg_13 ( .CK(CLK60M), .D(CRCREG199_13), .S(STSRST_), .Q(C13), 
        .QN(CRC[2]) );
    zdffsd CRCREG_reg_12 ( .CK(CLK60M), .D(CRCREG199_12), .S(STSRST_), .Q(C12), 
        .QN(CRC[3]) );
    zdffsd CRCREG_reg_11 ( .CK(CLK60M), .D(CRCREG199_11), .S(STSRST_), .Q(C11), 
        .QN(CRC[4]) );
    zdffsd CRCREG_reg_10 ( .CK(CLK60M), .D(CRCREG199_10), .S(STSRST_), .Q(C10), 
        .QN(CRC[5]) );
    zdffsd CRCREG_reg_9 ( .CK(CLK60M), .D(CRCREG199_9), .S(STSRST_), .Q(C9), 
        .QN(CRC[6]) );
    zdffqsd PKTCRC16_reg_15 ( .CK(CLK60M), .D(PKTCRC16298_15), .S(STSRST_), 
        .Q(PKTCRC16_15) );
    zdffqsd PKTCRC16_reg_9 ( .CK(CLK60M), .D(PKTCRC16298_9), .S(STSRST_), .Q(
        PKTCRC16_9) );
    zdffqsd PKTCRC16_reg_6 ( .CK(CLK60M), .D(PKTCRC16298_6), .S(STSRST_), .Q(
        PKTCRC16_6) );
    zdffqsd PKTCRC16_reg_5 ( .CK(CLK60M), .D(PKTCRC16298_5), .S(STSRST_), .Q(
        PKTCRC16_5) );
    zdffqsd PKTCRC16_reg_3 ( .CK(CLK60M), .D(PKTCRC16298_3), .S(STSRST_), .Q(
        PKTCRC16_3) );
    zao211b U265 ( .A(n411), .B(n415), .C(n409), .D(n416), .Y(CRCREG199_0) );
    zao211b U266 ( .A(n411), .B(n417), .C(n409), .D(n418), .Y(CRCREG199_1) );
    zao211b U267 ( .A(n411), .B(n419), .C(n409), .D(n420), .Y(CRCREG199_2) );
    zao211b U268 ( .A(n412), .B(n421), .C(n405), .D(n422), .Y(CRCREG199_3) );
    zao211b U269 ( .A(n412), .B(n423), .C(CRCRST), .D(n424), .Y(CRCREG199_4)
         );
    zao211b U270 ( .A(n412), .B(n425), .C(CRCRST), .D(n426), .Y(CRCREG199_5)
         );
    zao211b U271 ( .A(n412), .B(n427), .C(CRCRST), .D(n428), .Y(CRCREG199_6)
         );
    zao211b U272 ( .A(n411), .B(n429), .C(n405), .D(n430), .Y(CRCREG199_7) );
    zao211b U273 ( .A(n412), .B(n431), .C(n405), .D(n432), .Y(CRCREG199_8) );
    zao211b U274 ( .A(n411), .B(n433), .C(CRCRST), .D(n434), .Y(CRCREG199_9)
         );
    zao211b U275 ( .A(n548), .B(C10), .C(CRCRST), .D(n435), .Y(CRCREG199_10)
         );
    zao211b U276 ( .A(n_989), .B(n386), .C(n409), .D(n436), .Y(CRCREG199_11)
         );
    zao211b U277 ( .A(n_988), .B(n386), .C(n546), .D(n437), .Y(CRCREG199_12)
         );
    zao211b U278 ( .A(n_987), .B(n386), .C(n546), .D(n438), .Y(CRCREG199_13)
         );
    zao211b U279 ( .A(n_986), .B(n386), .C(n546), .D(n439), .Y(CRCREG199_14)
         );
    zao211b U280 ( .A(n_985), .B(n386), .C(n546), .D(n440), .Y(CRCREG199_15)
         );
    zao222b U281 ( .A(ADRENDPS[0]), .B(n546), .C(CRCHOLD_8), .D(n547), .E(n548
        ), .F(h0), .Y(CRCHOLD224_0) );
    zao222b U282 ( .A(ADRENDPS[1]), .B(n405), .C(CRCHOLD_9), .D(n412), .E(n407
        ), .F(h1), .Y(CRCHOLD224_1) );
    zao222b U283 ( .A(ADRENDPS[2]), .B(n409), .C(CRCHOLD_10), .D(n547), .E(
        n408), .F(h2), .Y(CRCHOLD224_2) );
    zao222b U284 ( .A(ADRENDPS[3]), .B(n405), .C(CRCHOLD_11), .D(n412), .E(
        n548), .F(h3), .Y(CRCHOLD224_3) );
    zao222b U285 ( .A(ADRENDPS[4]), .B(n409), .C(CRCHOLD_12), .D(n547), .E(
        n549), .F(h4), .Y(CRCHOLD224_4) );
    zao222b U286 ( .A(ADRENDPS[5]), .B(n405), .C(CRCHOLD_13), .D(n411), .E(
        n407), .F(h5), .Y(CRCHOLD224_5) );
    zao222b U287 ( .A(ADRENDPS[6]), .B(n405), .C(CRCHOLD_14), .D(n547), .E(
        n548), .F(h6), .Y(CRCHOLD224_6) );
    zao222b U288 ( .A(ADRENDPS[7]), .B(n409), .C(CRCHOLD_15), .D(n411), .E(
        n549), .F(h7), .Y(CRCHOLD224_7) );
    zao222b U289 ( .A(ADRENDPS[8]), .B(n405), .C(CRCHOLD_16), .D(n547), .E(
        CRCHOLD_8), .F(n549), .Y(CRCHOLD224_8) );
    zao222b U290 ( .A(n409), .B(ADRENDPS[9]), .C(CRCHOLD_17), .D(n547), .E(
        CRCHOLD_9), .F(n408), .Y(CRCHOLD224_9) );
    zao222b U291 ( .A(ADRENDPS[10]), .B(n405), .C(CRCHOLD_18), .D(n411), .E(
        CRCHOLD_10), .F(n548), .Y(CRCHOLD224_10) );
    zor2d U294 ( .A(n546), .B(n441), .Y(CRCSFT235_0) );
    zao211b U296 ( .A(PKTCRC16_0), .B(n407), .C(n409), .D(n442), .Y(
        PKTCRC16298_0) );
    zao211b U297 ( .A(PKTCRC16_1), .B(n408), .C(n546), .D(n443), .Y(
        PKTCRC16298_1) );
    zao211b U298 ( .A(PKTCRC16_2), .B(n548), .C(CRCRST), .D(n444), .Y(
        PKTCRC16298_2) );
    zao211b U299 ( .A(PKTCRC16_3), .B(n549), .C(n405), .D(n445), .Y(
        PKTCRC16298_3) );
    zao211b U300 ( .A(PKTCRC16_4), .B(n408), .C(n405), .D(n446), .Y(
        PKTCRC16298_4) );
    zao211b U301 ( .A(PKTCRC16_5), .B(n407), .C(n546), .D(n447), .Y(
        PKTCRC16298_5) );
    zao211b U302 ( .A(PKTCRC16_6), .B(n549), .C(CRCRST), .D(n448), .Y(
        PKTCRC16298_6) );
    zao211b U303 ( .A(PKTCRC16_7), .B(n408), .C(n546), .D(n449), .Y(
        PKTCRC16298_7) );
    zao211b U304 ( .A(PKTCRC16_8), .B(n548), .C(CRCRST), .D(n450), .Y(
        PKTCRC16298_8) );
    zao211b U305 ( .A(PKTCRC16_9), .B(n549), .C(n546), .D(n451), .Y(
        PKTCRC16298_9) );
    zao211b U306 ( .A(PKTCRC16_10), .B(n407), .C(n409), .D(n452), .Y(
        PKTCRC16298_10) );
    zao211b U307 ( .A(PKTCRC16_11), .B(n548), .C(n546), .D(n453), .Y(
        PKTCRC16298_11) );
    zao211b U308 ( .A(PKTCRC16_12), .B(n549), .C(n409), .D(n454), .Y(
        PKTCRC16298_12) );
    zao211b U309 ( .A(PKTCRC16_13), .B(n407), .C(n546), .D(n455), .Y(
        PKTCRC16298_13) );
    zao211b U310 ( .A(PKTCRC16_14), .B(n548), .C(n546), .D(n456), .Y(
        PKTCRC16298_14) );
    zao211b U311 ( .A(PKTCRC16_15), .B(n549), .C(n405), .D(n457), .Y(
        PKTCRC16298_15) );
    zan2d U312 ( .A(DATAIN[1]), .B(n411), .Y(n451) );
    zan2d U313 ( .A(DATAIN[0]), .B(n547), .Y(n450) );
    zan2d U314 ( .A(PKTCRC16_15), .B(n547), .Y(n449) );
    zan2d U315 ( .A(PKTCRC16_14), .B(n411), .Y(n448) );
    zan2d U316 ( .A(PKTCRC16_13), .B(n411), .Y(n447) );
    zan2d U317 ( .A(PKTCRC16_12), .B(n547), .Y(n446) );
    zan2d U318 ( .A(PKTCRC16_11), .B(n411), .Y(n445) );
    zan2d U319 ( .A(PKTCRC16_10), .B(n547), .Y(n444) );
    zan2d U320 ( .A(DATAIN[7]), .B(n411), .Y(n457) );
    zan2d U321 ( .A(DATAIN[6]), .B(n547), .Y(n456) );
    zan2d U322 ( .A(DATAIN[5]), .B(n547), .Y(n455) );
    zan2d U323 ( .A(DATAIN[4]), .B(n547), .Y(n454) );
    zan2d U324 ( .A(DATAIN[3]), .B(n547), .Y(n453) );
    zan2d U325 ( .A(DATAIN[2]), .B(n547), .Y(n452) );
    zan2d U326 ( .A(PKTCRC16_8), .B(n547), .Y(n442) );
    zan2d U327 ( .A(n549), .B(C9), .Y(n434) );
    zan2d U328 ( .A(n407), .B(CRCREG_6), .Y(n428) );
    zan2d U329 ( .A(n549), .B(CRCREG_3), .Y(n422) );
    zan2d U330 ( .A(n411), .B(CRCREG_2), .Y(n435) );
    zan2d U331 ( .A(n408), .B(CRCREG_0), .Y(n416) );
    zor2d U332 ( .A(n546), .B(n413), .Y(n463) );
    zivh U333 ( .A(DATAIN[2]), .Y(n475) );
    zxo2d U334 ( .A(C12), .B(n387), .Y(RC15) );
    zxo2d U335 ( .A(C11), .B(n388), .Y(RC14) );
    zxo2d U336 ( .A(n387), .B(n389), .Y(RC13) );
    zxo2d U337 ( .A(n389), .B(n482), .Y(RB15) );
    zxo2d U338 ( .A(n393), .B(n487), .Y(RB12) );
    zmux21ld U339 ( .A(n480), .B(n478), .S(n413), .Y(n441) );
    zor5b U340 ( .A(C15), .B(C11), .C(CRC[2]), .D(CRC[1]), .E(C12), .Y(n512)
         );
    zao211b U341 ( .A(MAC_SLAVE_ACT), .B(n514), .C(n515), .D(n516), .Y(n513)
         );
    zxo2d U342 ( .A(C12), .B(h3), .Y(n518) );
    zxo2d U343 ( .A(h5), .B(n518), .Y(n482) );
    zxo2d U344 ( .A(C12), .B(n390), .Y(n520) );
    zxo2d U345 ( .A(n392), .B(n520), .Y(n487) );
    zxo2d U346 ( .A(CRCREG_0), .B(n393), .Y(n490) );
    zxo2d U347 ( .A(C10), .B(C9), .Y(n522) );
    zxo2d U348 ( .A(DATAIN[5]), .B(n522), .Y(n493) );
    zxo2d U349 ( .A(CRCREG_7), .B(n393), .Y(n523) );
    zxo2d U350 ( .A(n399), .B(n402), .Y(n524) );
    zxo2d U351 ( .A(n403), .B(n524), .Y(n525) );
    zao22d U352 ( .A(n549), .B(C15), .C(n385), .D(n496), .Y(n440) );
    zao22d U353 ( .A(n549), .B(C14), .C(n385), .D(CRCREG_6), .Y(n439) );
    zao22d U354 ( .A(n548), .B(C13), .C(n385), .D(CRCREG_5), .Y(n438) );
    zao22d U355 ( .A(n549), .B(C12), .C(n385), .D(CRCREG_4), .Y(n437) );
    zao22d U356 ( .A(n549), .B(C11), .C(n385), .D(CRCREG_3), .Y(n436) );
    zxo2d U357 ( .A(C9), .B(DATAIN[6]), .Y(n526) );
    zxo2d U358 ( .A(C10), .B(n391), .Y(n530) );
    zxo2d U359 ( .A(DATAIN[1]), .B(n530), .Y(n531) );
    zxo2d U360 ( .A(n395), .B(n403), .Y(n532) );
    zxo2d U361 ( .A(n396), .B(n399), .Y(n502) );
    zor4b U362 ( .A(n506), .B(n507), .C(n504), .D(n505), .Y(n543) );
    zor4b U363 ( .A(CRCREG_7), .B(CRCREG_1), .C(C14), .D(C12), .Y(n544) );
    zor6b U364 ( .A(C10), .B(C9), .C(C11), .D(C13), .E(CRC[0]), .F(n544), .Y(
        n515) );
    zor4b U365 ( .A(CRCREG_4), .B(CRCREG_6), .C(CRCREG_5), .D(CRC[12]), .Y(
        n545) );
    zor4b U366 ( .A(CRCREG_8), .B(CRC[15]), .C(CRC[13]), .D(n545), .Y(n516) );
    zor6b U367 ( .A(n510), .B(n511), .C(n508), .D(n509), .E(n543), .F(n534), 
        .Y(n514) );
    zxo2d U368 ( .A(n475), .B(n395), .Y(n491) );
    zivh U369 ( .A(n464), .Y(n547) );
    zivh U370 ( .A(n463), .Y(n548) );
    zivh U371 ( .A(n463), .Y(n549) );
    zao22b U372 ( .A(CRCSFT_1), .B(n408), .C(CRCSFT_0), .D(n411), .Y(
        CRCSFT235_1) );
    zbfb U373 ( .A(CRCHOLD224_11), .Y(n550) );
    zbfb U374 ( .A(CRCHOLD224_12), .Y(n551) );
    zbfb U375 ( .A(CRCHOLD224_13), .Y(n552) );
    zao22b U376 ( .A(CRCHOLD_13), .B(n408), .C(ADRENDPS[13]), .D(n405), .Y(
        CRCHOLD224_13) );
    zbfb U377 ( .A(CRCHOLD224_14), .Y(n553) );
    zbfb U378 ( .A(CRCHOLD224_15), .Y(n554) );
    zbfb U379 ( .A(CRCHOLD224_16), .Y(n555) );
    zao22b U380 ( .A(CRCHOLD_16), .B(n407), .C(ADRENDPS[16]), .D(CRCRST), .Y(
        CRCHOLD224_16) );
    zbfb U381 ( .A(CRCHOLD224_17), .Y(n556) );
    zbfb U382 ( .A(CRCHOLD224_18), .Y(n557) );
endmodule


module MACETC ( MAC_ASKREPLY, ASKREPLY, EN_UTM_RESET, TXCRCEN, RXCRCEN, CRCEN, 
    TXCRCDAT, RXCRCDAT, CRCDATIN, TXCRCRST, RXCRCRST, CRCRST, DATPKT, RXDATA, 
    CRC16, TXADDR, TXENDP, SOFV, TXSOF, ADRENDPS, SPLIT, HUBADDR, SP_SC, 
    HUBPORT, SP_S, SP_E, SP_ET, NEWCMD, TRST_, STSRST_, HRST_, HCRESET, TXBCNT, 
    RXBCNT, ACTLEN, TD_IN, USBPOP, LIGHTRST, EHCIEXE, CLK60M, EOF1, EOF2, 
    T_EOF1, T_EOF2, CMDSTART, MAXLEN, SL_MAXLEN, MAC_MAXLEN, MAC_CMDSTART, 
    SLAVE_ACT, MAC_SLAVE_ACT, TXCRCPHASE, PTstCtrl_A_3, PTstCtrl_A_2, 
    PTstCtrl_A_1, PTstCtrl_A_0, PTstCtrl_B_3, PTstCtrl_B_2, PTstCtrl_B_1, 
    PTstCtrl_B_0, PTstCtrl_C_3, PTstCtrl_C_2, PTstCtrl_C_1, PTstCtrl_C_0, 
    PTstCtrl_D_3, PTstCtrl_D_2, PTstCtrl_D_1, PTstCtrl_D_0, PTstCtrl_E_3, 
    PTstCtrl_E_2, PTstCtrl_E_1, PTstCtrl_E_0, PTstCtrl_F_3, PTstCtrl_F_2, 
    PTstCtrl_F_1, PTstCtrl_F_0, PTstCtrl_G_3, PTstCtrl_G_2, PTstCtrl_G_1, 
    PTstCtrl_G_0, PTstCtrl_H_3, PTstCtrl_H_2, PTstCtrl_H_1, PTstCtrl_H_0, 
    PTEST_3, PTEST_2, PTEST_1, PTEST_0, TEST_J, TEST_K, TEST_PACKET, 
    TEST_FORCE_ENABLE, UTM_SOF, RXACTIVE, TXVALID, BABOPT, FBABBLE, 
    TEST_EYE_EN, TEST_EYE, ATPG_ENI, HS_TRST_, UTM_TXREADY, TXREADY_SYNC, 
    UTM_RUN );
input  [7:0] TXCRCDAT;
input  [7:0] RXCRCDAT;
input  [3:0] TXENDP;
input  [6:0] HUBPORT;
input  [6:0] TXADDR;
output [18:0] ADRENDPS;
input  [6:0] HUBADDR;
input  [1:0] SP_ET;
output [10:0] MAC_MAXLEN;
output [7:0] CRCDATIN;
input  [10:0] SOFV;
output [10:0] ACTLEN;
input  [10:0] SL_MAXLEN;
input  [10:0] TXBCNT;
input  [10:0] RXBCNT;
input  [10:0] MAXLEN;
input  MAC_ASKREPLY, EN_UTM_RESET, TXCRCEN, RXCRCEN, TXCRCRST, RXCRCRST, 
    DATPKT, RXDATA, TXSOF, SPLIT, SP_SC, SP_S, SP_E, NEWCMD, HRST_, HCRESET, 
    TD_IN, USBPOP, LIGHTRST, EHCIEXE, CLK60M, EOF1, EOF2, CMDSTART, SLAVE_ACT, 
    TXCRCPHASE, PTstCtrl_A_3, PTstCtrl_A_2, PTstCtrl_A_1, PTstCtrl_A_0, 
    PTstCtrl_B_3, PTstCtrl_B_2, PTstCtrl_B_1, PTstCtrl_B_0, PTstCtrl_C_3, 
    PTstCtrl_C_2, PTstCtrl_C_1, PTstCtrl_C_0, PTstCtrl_D_3, PTstCtrl_D_2, 
    PTstCtrl_D_1, PTstCtrl_D_0, PTstCtrl_E_3, PTstCtrl_E_2, PTstCtrl_E_1, 
    PTstCtrl_E_0, PTstCtrl_F_3, PTstCtrl_F_2, PTstCtrl_F_1, PTstCtrl_F_0, 
    PTstCtrl_G_3, PTstCtrl_G_2, PTstCtrl_G_1, PTstCtrl_G_0, PTstCtrl_H_3, 
    PTstCtrl_H_2, PTstCtrl_H_1, PTstCtrl_H_0, RXACTIVE, TXVALID, BABOPT, 
    TEST_EYE_EN, ATPG_ENI, HS_TRST_, UTM_TXREADY, UTM_RUN;
output ASKREPLY, CRCEN, CRCRST, CRC16, TRST_, STSRST_, T_EOF1, T_EOF2, 
    MAC_CMDSTART, MAC_SLAVE_ACT, PTEST_3, PTEST_2, PTEST_1, PTEST_0, TEST_J, 
    TEST_K, TEST_PACKET, TEST_FORCE_ENABLE, UTM_SOF, FBABBLE, TEST_EYE, 
    TXREADY_SYNC;
    wire ACTLEN911_7, SPAREO6, TESTM_T1093, TESTM_T, UTM_SOF_T, SPAREO0_, 
        SPAREO8, ACTLEN911_10, UTM_SOF_T1185, ACTLEN911_9, SPAREO1, 
        ACTLEN911_0, ACTLEN911_8, SPAREO9, ACTLEN911_1, SPAREO0, SPAREO7, 
        ACTLEN911_6, STSRST_PRE, TESTM_2T, STSRST_PRE835, ACTLEN911_4, SPAREO5, 
        TESTM_3T, UTM_SOF_2T, SPAREO2, ACTLEN911_3, ACTLEN911_2, SPAREO3, 
        SPAREO1_, EHCIEXE_T, EHCIEXE_2T, SPAREO4, ACTLEN911_5, n1299, n1300, 
        n1301, n1302, n1303, n1304, n1305, n1307, n1316, n1317, n1318, n1319, 
        n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
        n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
        n1340, n1341, n1342, n1343, n1344, n1345;
    zaoi211b SPARE672 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE675 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zoai21b SPARE674 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE673 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zivb SPARE678 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE671 ( .CK(CLK60M), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    znr3b SPARE676 ( .A(SPAREO2), .B(EHCIEXE_2T), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE677 ( .A(SPAREO4), .Y(SPAREO5) );
    znd3b SPARE679 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE670 ( .CK(CLK60M), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znr2b U263 ( .A(HCRESET), .B(LIGHTRST), .Y(n1323) );
    zor2b U264 ( .A(n1330), .B(TXSOF), .Y(UTM_SOF_T1185) );
    zivb U265 ( .A(TD_IN), .Y(n1338) );
    znr2b U266 ( .A(NEWCMD), .B(n1326), .Y(STSRST_PRE835) );
    zan3b U267 ( .A(n1325), .B(TEST_EYE_EN), .C(TESTM_3T), .Y(TEST_EYE) );
    zivb U268 ( .A(n1328), .Y(n1325) );
    zivb U269 ( .A(n1332), .Y(n1336) );
    zcx4b U270 ( .A(RXACTIVE), .B(TXVALID), .C(n1318), .D(BABOPT), .Y(FBABBLE)
         );
    zor2b U271 ( .A(n1324), .B(UTM_RUN), .Y(UTM_SOF) );
    zan3b U272 ( .A(n1305), .B(PTEST_2), .C(TESTM_3T), .Y(TEST_FORCE_ENABLE)
         );
    zan3b U273 ( .A(n1304), .B(n1317), .C(TESTM_3T), .Y(TEST_K) );
    zan3b U274 ( .A(n1305), .B(n1319), .C(TESTM_3T), .Y(TEST_J) );
    zivb U275 ( .A(PTEST_0), .Y(n1317) );
    zivb U276 ( .A(PTEST_1), .Y(n1335) );
    zivb U277 ( .A(PTEST_2), .Y(n1319) );
    zmux21hb U278 ( .A(MAXLEN[0]), .B(SL_MAXLEN[0]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[0]) );
    zmux21hb U279 ( .A(MAXLEN[1]), .B(SL_MAXLEN[1]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[1]) );
    zmux21hb U280 ( .A(MAXLEN[2]), .B(SL_MAXLEN[2]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[2]) );
    zmux21hb U281 ( .A(MAXLEN[3]), .B(SL_MAXLEN[3]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[3]) );
    zmux21hb U282 ( .A(MAXLEN[4]), .B(SL_MAXLEN[4]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[4]) );
    zmux21hb U283 ( .A(MAXLEN[5]), .B(SL_MAXLEN[5]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[5]) );
    zmux21hb U284 ( .A(MAXLEN[6]), .B(SL_MAXLEN[6]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[6]) );
    zmux21hb U285 ( .A(MAXLEN[7]), .B(SL_MAXLEN[7]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[7]) );
    zmux21hb U286 ( .A(MAXLEN[8]), .B(SL_MAXLEN[8]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[8]) );
    zmux21hb U287 ( .A(MAXLEN[9]), .B(SL_MAXLEN[9]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[9]) );
    zmux21hb U288 ( .A(MAXLEN[10]), .B(SL_MAXLEN[10]), .S(MAC_SLAVE_ACT), .Y(
        MAC_MAXLEN[10]) );
    zivb U289 ( .A(n1318), .Y(T_EOF2) );
    zivb U290 ( .A(EOF2), .Y(n1334) );
    zan3b U291 ( .A(EOF1), .B(n1321), .C(n1322), .Y(T_EOF1) );
    zor2b U292 ( .A(n1332), .B(n1333), .Y(n1322) );
    zivb U293 ( .A(n1322), .Y(TEST_PACKET) );
    zivb U294 ( .A(SPLIT), .Y(n1337) );
    zmux21hb U295 ( .A(DATPKT), .B(RXDATA), .S(MAC_ASKREPLY), .Y(CRC16) );
    zmux21hb U296 ( .A(TXCRCRST), .B(RXCRCRST), .S(MAC_ASKREPLY), .Y(CRCRST)
         );
    zmux21hb U297 ( .A(TXCRCDAT[0]), .B(RXCRCDAT[0]), .S(MAC_ASKREPLY), .Y(
        CRCDATIN[0]) );
    zmux21hb U298 ( .A(TXCRCDAT[1]), .B(RXCRCDAT[1]), .S(MAC_ASKREPLY), .Y(
        CRCDATIN[1]) );
    zmux21hb U299 ( .A(TXCRCDAT[2]), .B(RXCRCDAT[2]), .S(MAC_ASKREPLY), .Y(
        CRCDATIN[2]) );
    zmux21hb U300 ( .A(TXCRCDAT[3]), .B(RXCRCDAT[3]), .S(MAC_ASKREPLY), .Y(
        CRCDATIN[3]) );
    zmux21hb U301 ( .A(TXCRCDAT[4]), .B(RXCRCDAT[4]), .S(MAC_ASKREPLY), .Y(
        CRCDATIN[4]) );
    zmux21hb U302 ( .A(TXCRCDAT[5]), .B(RXCRCDAT[5]), .S(MAC_ASKREPLY), .Y(
        CRCDATIN[5]) );
    zmux21hb U303 ( .A(TXCRCDAT[6]), .B(RXCRCDAT[6]), .S(MAC_ASKREPLY), .Y(
        CRCDATIN[6]) );
    zmux21hb U304 ( .A(TXCRCDAT[7]), .B(RXCRCDAT[7]), .S(MAC_ASKREPLY), .Y(
        CRCDATIN[7]) );
    zaoi21b U305 ( .A(EN_UTM_RESET), .B(EOF2), .C(n1331), .Y(ASKREPLY) );
    zivb U306 ( .A(MAC_ASKREPLY), .Y(n1331) );
    zivb U307 ( .A(TESTM_3T), .Y(n1333) );
    zivb U308 ( .A(MAC_SLAVE_ACT), .Y(n1321) );
    znr2b U309 ( .A(TXCRCPHASE), .B(CRCEN), .Y(n1299) );
    znr2b U310 ( .A(TXSOF), .B(n1337), .Y(n1300) );
    znr2b U311 ( .A(TXSOF), .B(SPLIT), .Y(n1301) );
    znr2b U312 ( .A(n1299), .B(n1338), .Y(n1302) );
    znr2b U313 ( .A(n1299), .B(TD_IN), .Y(n1303) );
    znr3b U314 ( .A(PTEST_2), .B(PTEST_3), .C(n1335), .Y(n1304) );
    znr3b U315 ( .A(PTEST_1), .B(PTEST_3), .C(n1317), .Y(n1305) );
    zmux21hb U316 ( .A(TXCRCEN), .B(RXCRCEN), .S(MAC_ASKREPLY), .Y(CRCEN) );
    zbfb U317 ( .A(HS_TRST_), .Y(n1307) );
    zdffqrb_ MAC_SLAVE_ACT_reg ( .CK(CLK60M), .D(SLAVE_ACT), .R(n1307), .Q(
        MAC_SLAVE_ACT) );
    zdffqrb_ MAC_CMDSTART_reg ( .CK(CLK60M), .D(CMDSTART), .R(n1307), .Q(
        MAC_CMDSTART) );
    zdffqrb TESTM_T_reg ( .CK(CLK60M), .D(TESTM_T1093), .R(HS_TRST_), .Q(
        TESTM_T) );
    zdffqrb EHCIEXE_T_reg ( .CK(CLK60M), .D(EHCIEXE), .R(n1307), .Q(EHCIEXE_T)
         );
    zdffqrb TESTM_2T_reg ( .CK(CLK60M), .D(n1345), .R(n1307), .Q(TESTM_2T) );
    zdffqrb STSRST_PRE_reg ( .CK(CLK60M), .D(STSRST_PRE835), .R(n1307), .Q(
        STSRST_PRE) );
    zdffqrb TXREADY_SYNC_reg ( .CK(CLK60M), .D(UTM_TXREADY), .R(n1307), .Q(
        TXREADY_SYNC) );
    zdffqrb EHCIEXE_2T_reg ( .CK(CLK60M), .D(n1343), .R(n1307), .Q(EHCIEXE_2T)
         );
    zdffqrb_ UTM_SOF_2T_reg ( .CK(CLK60M), .D(n1339), .R(HS_TRST_), .Q(
        UTM_SOF_2T) );
    zdffqrb_ ACTLEN_reg_0 ( .CK(CLK60M), .D(ACTLEN911_0), .R(HS_TRST_), .Q(
        ACTLEN[0]) );
    zdffqrb_ ACTLEN_reg_3 ( .CK(CLK60M), .D(ACTLEN911_3), .R(HS_TRST_), .Q(
        ACTLEN[3]) );
    zdffqrb_ ACTLEN_reg_9 ( .CK(CLK60M), .D(ACTLEN911_9), .R(HS_TRST_), .Q(
        ACTLEN[9]) );
    zdffqrb_ ACTLEN_reg_8 ( .CK(CLK60M), .D(ACTLEN911_8), .R(HS_TRST_), .Q(
        ACTLEN[8]) );
    zdffqrb_ ACTLEN_reg_4 ( .CK(CLK60M), .D(ACTLEN911_4), .R(HS_TRST_), .Q(
        ACTLEN[4]) );
    zdffqrb_ TESTM_3T_reg ( .CK(CLK60M), .D(TESTM_2T), .R(HS_TRST_), .Q(
        TESTM_3T) );
    zdffqrb_ ACTLEN_reg_10 ( .CK(CLK60M), .D(ACTLEN911_10), .R(HS_TRST_), .Q(
        ACTLEN[10]) );
    zdffqrb_ ACTLEN_reg_1 ( .CK(CLK60M), .D(ACTLEN911_1), .R(HS_TRST_), .Q(
        ACTLEN[1]) );
    zdffqrb_ UTM_SOF_T_reg ( .CK(CLK60M), .D(UTM_SOF_T1185), .R(HS_TRST_), .Q(
        UTM_SOF_T) );
    zdffqrb_ ACTLEN_reg_5 ( .CK(CLK60M), .D(ACTLEN911_5), .R(HS_TRST_), .Q(
        ACTLEN[5]) );
    zdffqrb_ ACTLEN_reg_2 ( .CK(CLK60M), .D(ACTLEN911_2), .R(HS_TRST_), .Q(
        ACTLEN[2]) );
    zdffqrb_ ACTLEN_reg_6 ( .CK(CLK60M), .D(ACTLEN911_6), .R(HS_TRST_), .Q(
        ACTLEN[6]) );
    zdffqrb_ ACTLEN_reg_7 ( .CK(CLK60M), .D(ACTLEN911_7), .R(HS_TRST_), .Q(
        ACTLEN[7]) );
    zbfb U318 ( .A(HUBPORT[3]), .Y(ADRENDPS[11]) );
    zbfb U319 ( .A(HUBPORT[4]), .Y(ADRENDPS[12]) );
    zbfb U320 ( .A(HUBPORT[5]), .Y(ADRENDPS[13]) );
    zbfb U321 ( .A(HUBPORT[6]), .Y(ADRENDPS[14]) );
    zbfb U322 ( .A(SP_S), .Y(ADRENDPS[15]) );
    zbfb U323 ( .A(SP_E), .Y(ADRENDPS[16]) );
    zbfb U324 ( .A(SP_ET[0]), .Y(ADRENDPS[17]) );
    zbfb U325 ( .A(SP_ET[1]), .Y(ADRENDPS[18]) );
    zor5b U326 ( .A(PTstCtrl_A_2), .B(PTstCtrl_B_2), .C(PTstCtrl_E_2), .D(
        PTstCtrl_C_2), .E(n1316), .Y(PTEST_2) );
    zor5b U327 ( .A(PTstCtrl_F_0), .B(PTstCtrl_E_0), .C(PTstCtrl_A_0), .D(
        PTstCtrl_B_0), .E(n1320), .Y(PTEST_0) );
    zao21d U328 ( .A(n1323), .B(HRST_), .C(ATPG_ENI), .Y(TRST_) );
    zor5b U329 ( .A(PTstCtrl_G_1), .B(PTstCtrl_E_1), .C(PTstCtrl_B_1), .D(
        PTstCtrl_D_1), .E(n1327), .Y(PTEST_1) );
    zor3b U330 ( .A(TEST_EYE_EN), .B(n1304), .C(n1328), .Y(TESTM_T1093) );
    zor2d U331 ( .A(STSRST_PRE), .B(ATPG_ENI), .Y(STSRST_) );
    zor5b U332 ( .A(PTstCtrl_B_3), .B(PTstCtrl_E_3), .C(PTstCtrl_D_3), .D(
        PTstCtrl_C_3), .E(n1329), .Y(PTEST_3) );
    zao222b U333 ( .A(RXBCNT[10]), .B(n1302), .C(TXBCNT[10]), .D(n1303), .E(
        ACTLEN[10]), .F(n1299), .Y(ACTLEN911_10) );
    zao222b U334 ( .A(RXBCNT[9]), .B(n1302), .C(TXBCNT[9]), .D(n1303), .E(
        n1299), .F(ACTLEN[9]), .Y(ACTLEN911_9) );
    zao222b U335 ( .A(RXBCNT[8]), .B(n1302), .C(TXBCNT[8]), .D(n1303), .E(
        ACTLEN[8]), .F(n1299), .Y(ACTLEN911_8) );
    zao222b U336 ( .A(RXBCNT[7]), .B(n1302), .C(TXBCNT[7]), .D(n1303), .E(
        ACTLEN[7]), .F(n1299), .Y(ACTLEN911_7) );
    zao222b U337 ( .A(RXBCNT[6]), .B(n1302), .C(TXBCNT[6]), .D(n1303), .E(
        ACTLEN[6]), .F(n1299), .Y(ACTLEN911_6) );
    zao222b U338 ( .A(RXBCNT[5]), .B(n1302), .C(TXBCNT[5]), .D(n1303), .E(
        ACTLEN[5]), .F(n1299), .Y(ACTLEN911_5) );
    zao222b U339 ( .A(RXBCNT[4]), .B(n1302), .C(TXBCNT[4]), .D(n1303), .E(
        ACTLEN[4]), .F(n1299), .Y(ACTLEN911_4) );
    zao222b U340 ( .A(RXBCNT[3]), .B(n1302), .C(TXBCNT[3]), .D(n1303), .E(
        ACTLEN[3]), .F(n1299), .Y(ACTLEN911_3) );
    zao222b U341 ( .A(RXBCNT[2]), .B(n1302), .C(TXBCNT[2]), .D(n1303), .E(
        ACTLEN[2]), .F(n1299), .Y(ACTLEN911_2) );
    zao222b U342 ( .A(RXBCNT[1]), .B(n1302), .C(TXBCNT[1]), .D(n1303), .E(
        ACTLEN[1]), .F(n1299), .Y(ACTLEN911_1) );
    zao222b U343 ( .A(RXBCNT[0]), .B(n1302), .C(TXBCNT[0]), .D(n1303), .E(
        ACTLEN[0]), .F(n1299), .Y(ACTLEN911_0) );
    zao222b U344 ( .A(HUBPORT[2]), .B(n1300), .C(TXENDP[3]), .D(n1301), .E(
        SOFV[10]), .F(TXSOF), .Y(ADRENDPS[10]) );
    zao222b U345 ( .A(HUBPORT[1]), .B(n1300), .C(TXENDP[2]), .D(n1301), .E(
        TXSOF), .F(SOFV[9]), .Y(ADRENDPS[9]) );
    zao222b U346 ( .A(HUBPORT[0]), .B(n1300), .C(TXENDP[1]), .D(n1301), .E(
        SOFV[8]), .F(TXSOF), .Y(ADRENDPS[8]) );
    zao222b U347 ( .A(SP_SC), .B(n1300), .C(TXENDP[0]), .D(n1301), .E(SOFV[7]), 
        .F(TXSOF), .Y(ADRENDPS[7]) );
    zao222b U348 ( .A(HUBADDR[6]), .B(n1300), .C(TXADDR[6]), .D(n1301), .E(
        SOFV[6]), .F(TXSOF), .Y(ADRENDPS[6]) );
    zao222b U349 ( .A(HUBADDR[5]), .B(n1300), .C(TXADDR[5]), .D(n1301), .E(
        SOFV[5]), .F(TXSOF), .Y(ADRENDPS[5]) );
    zao222b U350 ( .A(HUBADDR[4]), .B(n1300), .C(TXADDR[4]), .D(n1301), .E(
        SOFV[4]), .F(TXSOF), .Y(ADRENDPS[4]) );
    zao222b U351 ( .A(HUBADDR[3]), .B(n1300), .C(TXADDR[3]), .D(n1301), .E(
        SOFV[3]), .F(TXSOF), .Y(ADRENDPS[3]) );
    zao222b U352 ( .A(HUBADDR[2]), .B(n1300), .C(TXADDR[2]), .D(n1301), .E(
        SOFV[2]), .F(TXSOF), .Y(ADRENDPS[2]) );
    zao222b U353 ( .A(HUBADDR[1]), .B(n1300), .C(TXADDR[1]), .D(n1301), .E(
        SOFV[1]), .F(TXSOF), .Y(ADRENDPS[1]) );
    zao222b U354 ( .A(HUBADDR[0]), .B(n1300), .C(TXADDR[0]), .D(n1301), .E(
        SOFV[0]), .F(TXSOF), .Y(ADRENDPS[0]) );
    zinr2b U355 ( .A(TESTM_T), .B(TESTM_2T), .Y(n1330) );
    zinr2b U356 ( .A(UTM_SOF_T), .B(UTM_SOF_2T), .Y(n1324) );
    zinr2b U357 ( .A(EHCIEXE_T), .B(EHCIEXE_2T), .Y(n1326) );
    zor4b U358 ( .A(PTEST_3), .B(n1319), .C(PTEST_0), .D(PTEST_1), .Y(n1332)
         );
    zao211b U359 ( .A(n1304), .B(n1317), .C(n1336), .D(n1305), .Y(n1328) );
    zor3b U360 ( .A(MAC_SLAVE_ACT), .B(n1334), .C(TEST_PACKET), .Y(n1318) );
    zor4b U361 ( .A(PTstCtrl_G_0), .B(PTstCtrl_D_0), .C(PTstCtrl_H_0), .D(
        PTstCtrl_C_0), .Y(n1320) );
    zor4b U362 ( .A(PTstCtrl_H_1), .B(PTstCtrl_F_1), .C(PTstCtrl_A_1), .D(
        PTstCtrl_C_1), .Y(n1327) );
    zor4b U363 ( .A(PTstCtrl_A_3), .B(PTstCtrl_H_3), .C(PTstCtrl_G_3), .D(
        PTstCtrl_F_3), .Y(n1329) );
    zor4b U364 ( .A(PTstCtrl_G_2), .B(PTstCtrl_F_2), .C(PTstCtrl_H_2), .D(
        PTstCtrl_D_2), .Y(n1316) );
    zbfb U365 ( .A(n1341), .Y(n1339) );
    zivb U366 ( .A(UTM_SOF_T), .Y(n1340) );
    zivb U367 ( .A(n1340), .Y(n1341) );
    zivb U368 ( .A(EHCIEXE_T), .Y(n1342) );
    zivb U369 ( .A(n1342), .Y(n1343) );
    zivb U370 ( .A(TESTM_T), .Y(n1344) );
    zivb U371 ( .A(n1344), .Y(n1345) );
endmodule


module HS_PIDENC ( TXOUT, TXIN, TXSOF, TXSETUP, TXDATA0, TXDATA1, TXDATA2, 
    TXMDATA, TXACK, TXNAK, TXSTALL, TXNYET, TXERR, TXSPLIT, TXPING, TX_PID, 
    TOKEN, DATPKT, HANDSHK, SPLIT, MAC_SLAVE_ACT, SL_PID, SL_FORCE_PID );
output [7:0] TX_PID;
input  [3:0] SL_PID;
input  TXOUT, TXIN, TXSOF, TXSETUP, TXDATA0, TXDATA1, TXDATA2, TXMDATA, TXACK, 
    TXNAK, TXSTALL, TXNYET, TXERR, TXSPLIT, TXPING, MAC_SLAVE_ACT, 
    SL_FORCE_PID;
output TOKEN, DATPKT, HANDSHK, SPLIT;
    wire n498, n499, n500, n501, n502, n503, n504, n505, n506;
    zbfb U99 ( .A(TXSPLIT), .Y(SPLIT) );
    zao22b U100 ( .A(MAC_SLAVE_ACT), .B(SL_PID[3]), .C(n498), .D(n499), .Y(
        TX_PID[3]) );
    zao22b U101 ( .A(SL_PID[2]), .B(MAC_SLAVE_ACT), .C(n498), .D(n500), .Y(
        TX_PID[2]) );
    zor4b U102 ( .A(TXDATA0), .B(TXMDATA), .C(TXDATA2), .D(TXDATA1), .Y(DATPKT
        ) );
    zor2b U103 ( .A(TXERR), .B(n501), .Y(HANDSHK) );
    zor3b U104 ( .A(TXPING), .B(TXSPLIT), .C(n502), .Y(TOKEN) );
    znr4b U105 ( .A(TXNYET), .B(TXPING), .C(TXSOF), .D(TXDATA2), .Y(n499) );
    znr4b U106 ( .A(TXOUT), .B(TXACK), .C(MAC_SLAVE_ACT), .D(TXDATA0), .Y(n498
        ) );
    zor4b U107 ( .A(TXACK), .B(TXSTALL), .C(TXNYET), .D(TXNAK), .Y(n501) );
    zor4b U108 ( .A(TXOUT), .B(TXSETUP), .C(TXSOF), .D(TXIN), .Y(n502) );
    zxn2b U109 ( .A(SL_FORCE_PID), .B(TX_PID[3]), .Y(TX_PID[7]) );
    zxn2b U110 ( .A(SL_FORCE_PID), .B(TX_PID[2]), .Y(TX_PID[6]) );
    zoa21b U111 ( .A(DATPKT), .B(n501), .C(n504), .Y(n503) );
    zor2b U112 ( .A(n502), .B(DATPKT), .Y(n505) );
    zxn2b U113 ( .A(TX_PID[1]), .B(SL_FORCE_PID), .Y(TX_PID[5]) );
    zxn2b U114 ( .A(TX_PID[0]), .B(SL_FORCE_PID), .Y(TX_PID[4]) );
    zor4b U115 ( .A(TXNAK), .B(TXSPLIT), .C(TXIN), .D(TXDATA1), .Y(n506) );
    znd2b U116 ( .A(n499), .B(n506), .Y(n500) );
    zivb U117 ( .A(n502), .Y(n504) );
    zmux21hb U118 ( .A(n503), .B(SL_PID[1]), .S(MAC_SLAVE_ACT), .Y(TX_PID[1])
         );
    zmux21hb U119 ( .A(n505), .B(SL_PID[0]), .S(MAC_SLAVE_ACT), .Y(TX_PID[0])
         );
endmodule


module HS_PIDEC ( RXPID, RXACK, RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXDATA, 
    RXNAK, RXSTALL, RXNYET, RXERR, RXHAND, RXTOKEN, PIDERR, RXOUT, RXIN, RXSOF, 
    RXSETUP, RXPING, RXSPLIT, LATCHPID, STSRST_, ISO, SEQERR, MAC_SLAVE_ACT, 
    ENISOHANDCHK, ATPG_ENI );
input  [7:0] RXPID;
input  LATCHPID, STSRST_, ISO, SEQERR, MAC_SLAVE_ACT, ENISOHANDCHK, ATPG_ENI;
output RXACK, RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXDATA, RXNAK, RXSTALL, 
    RXNYET, RXERR, RXHAND, RXTOKEN, PIDERR, RXOUT, RXIN, RXSOF, RXSETUP, 
    RXPING, RXSPLIT;
    wire val228_1, n208, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
        n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
        n305;
    zlthqrb PIDERR_reg ( .CK(n208), .D(val228_1), .R(STSRST_), .Q(PIDERR) );
    zor2b U109 ( .A(ATPG_ENI), .B(LATCHPID), .Y(n208) );
    zor3b U110 ( .A(SEQERR), .B(n284), .C(n285), .Y(val228_1) );
    zan2b U111 ( .A(n286), .B(n287), .Y(RXERR) );
    zan2b U112 ( .A(n288), .B(n289), .Y(RXNYET) );
    zan2b U113 ( .A(n287), .B(n290), .Y(RXSPLIT) );
    zan2b U114 ( .A(n287), .B(n288), .Y(RXPING) );
    zan2b U115 ( .A(n286), .B(n291), .Y(RXSETUP) );
    zan2b U116 ( .A(n291), .B(n288), .Y(RXSOF) );
    zan2b U117 ( .A(n291), .B(n292), .Y(RXOUT) );
    zan2b U118 ( .A(n290), .B(n291), .Y(RXIN) );
    zan2b U119 ( .A(n292), .B(n289), .Y(RXACK) );
    zan2b U120 ( .A(RXDATA), .B(n286), .Y(RXMDATA) );
    zan2b U121 ( .A(RXDATA), .B(n288), .Y(RXDATA2) );
    zan2b U122 ( .A(RXDATA), .B(n290), .Y(RXDATA1) );
    zan2b U123 ( .A(RXDATA), .B(n292), .Y(RXDATA0) );
    zan3b U124 ( .A(n289), .B(n293), .C(n290), .Y(RXNAK) );
    zan3b U125 ( .A(n286), .B(n293), .C(n289), .Y(RXSTALL) );
    znr3b U126 ( .A(n290), .B(RXPID[0]), .C(n288), .Y(n294) );
    zaoi21b U127 ( .A(n295), .B(n296), .C(MAC_SLAVE_ACT), .Y(n284) );
    zxo2b U128 ( .A(n298), .B(RXPID[5]), .Y(n297) );
    zxo2b U129 ( .A(n300), .B(RXPID[4]), .Y(n299) );
    zxo2b U130 ( .A(n302), .B(RXPID[7]), .Y(n301) );
    zxo2b U131 ( .A(n304), .B(RXPID[6]), .Y(n303) );
    zivb U132 ( .A(RXPID[1]), .Y(n298) );
    zivb U133 ( .A(RXPID[0]), .Y(n300) );
    zivb U134 ( .A(RXPID[3]), .Y(n302) );
    zivb U135 ( .A(RXPID[2]), .Y(n304) );
    zor4b U136 ( .A(n301), .B(n303), .C(n297), .D(n299), .Y(n285) );
    zcx4b U137 ( .A(RXPID[1]), .B(n286), .C(RXPID[0]), .D(n285), .Y(RXHAND) );
    zor2b U138 ( .A(n285), .B(RXPID[1]), .Y(n305) );
    zan2b U139 ( .A(RXPID[2]), .B(RXPID[3]), .Y(n286) );
    znr3b U140 ( .A(RXPID[0]), .B(n298), .C(n285), .Y(n289) );
    znr2b U141 ( .A(RXPID[0]), .B(n305), .Y(n287) );
    zan2b U142 ( .A(RXPID[3]), .B(n304), .Y(n290) );
    znr2b U143 ( .A(n300), .B(n305), .Y(n291) );
    zan2b U144 ( .A(RXPID[2]), .B(n302), .Y(n288) );
    zan2b U145 ( .A(n304), .B(n302), .Y(n292) );
    znr3b U146 ( .A(n298), .B(n300), .C(n285), .Y(RXDATA) );
    zor2b U147 ( .A(n294), .B(n305), .Y(n295) );
    zivb U148 ( .A(n295), .Y(RXTOKEN) );
    zivb U149 ( .A(PIDERR), .Y(n293) );
    znd3b U150 ( .A(RXHAND), .B(ENISOHANDCHK), .C(ISO), .Y(n296) );
endmodule


module HS_MACCTL ( NEWCMD, EOF1, EOF2, TD_IN, TD_OUT, TD_SETUP, TD_SPLIT, 
    TD_PING, MAC_CMDSTART, SOFGEN, CLK60M, ASKREPLY, ISO, TXSPLIT, TXACK, 
    TXDATA0, TXDATA1, TXDATA2, TXMDATA, TXIN, TXOUT, TXSOF, TXSETUP, TXPING, 
    TRST_, TXSTART, PKTXEND, PKRVEND, RXDATA, NORMPKT, SEQERR, W4REPLY, RXACK, 
    MAC_EOT, EOFTERM, DAT0, DAT1, DAT2, DATM, SP_SC, TEST_PACKET, 
    MAC_SLAVE_ACT, RXSOF, RXIN, RXOUT, RXSETUP, RXSPLIT, RXPING, RXTOKENPHASE, 
    DATAIN, PERIOD_CMD, ASYNC_CMD, RXADDRF, SL_PID, SL_TOGMATCH, RXPID, 
    SL_CRC16, SL_PERIOD, SL_DATA_PIDERR, SL_ET_ERR, SL_SE_ERR, SL_ACK_ERR, 
    SL_TXDATASEL, SL_TXFIXDATA, SL_MAXLEN, SL_FORCE_CRC, SL_FORCE_PID, 
    SL_FORCE_STUFF, DISPDRCV, RCV_POWERUP, TXTMOUT_EN, TMOUT_PARM, TXDELAY_EN, 
    TXDELAY_PARM, TURNCNT_EN, TX_PERIOD );
input  [31:0] PERIOD_CMD;
input  [23:0] RXADDRF;
input  [7:0] RXPID;
output [2:0] SL_TXDATASEL;
output [10:0] SL_MAXLEN;
output [7:0] SL_TXFIXDATA;
input  [7:0] TXDELAY_PARM;
input  [31:0] ASYNC_CMD;
output [3:0] SL_PID;
output [15:0] SL_CRC16;
input  [7:0] TMOUT_PARM;
input  EOF1, EOF2, TD_IN, TD_OUT, TD_SETUP, TD_SPLIT, TD_PING, MAC_CMDSTART, 
    SOFGEN, CLK60M, ISO, TRST_, PKTXEND, PKRVEND, RXDATA, NORMPKT, RXACK, DAT0, 
    DAT1, DAT2, DATM, SP_SC, TEST_PACKET, MAC_SLAVE_ACT, RXSOF, RXIN, RXOUT, 
    RXSETUP, RXSPLIT, RXPING, DISPDRCV, TXTMOUT_EN, TXDELAY_EN, TURNCNT_EN;
output NEWCMD, ASKREPLY, TXSPLIT, TXACK, TXDATA0, TXDATA1, TXDATA2, TXMDATA, 
    TXIN, TXOUT, TXSOF, TXSETUP, TXPING, TXSTART, SEQERR, W4REPLY, MAC_EOT, 
    EOFTERM, RXTOKENPHASE, DATAIN, SL_TOGMATCH, SL_PERIOD, SL_DATA_PIDERR, 
    SL_ET_ERR, SL_SE_ERR, SL_ACK_ERR, SL_FORCE_CRC, SL_FORCE_PID, 
    SL_FORCE_STUFF, RCV_POWERUP, TX_PERIOD;
    wire CMDSTATE_15, SL_RXSPLIT2598, SL_SP_ET2642_0, CMDSTATE_5, SPAREO6, 
        n2478, TXTMCNT2304_1, SL_DATA_PIDERR2868, TXDLCNT_5, TXTMCNT_1, 
        CMDSMNXT_14, TXTMCNT2296_2, CMDSMNXT_13, CMDSMNXT_5, TXDLCNT2426_7, 
        CMDSMNXT_2, TXDLCNT2418_0, TXDLCNT2418_7, SL_SP_S, EOFTERM2247, 
        TXDLCNT2426_0, SL_SP_ET_1, SPAREO0_, TXTMCNT2296_5, SPAREO8, W4SOFGEN, 
        TXTMCNT_6, TXTMCNT2304_6, TXDLCNT_2, SL_SE_ERR2808, SL_SP_E, 
        CMDSTATE_14, SPAREO1, CURISTX, TXTMCNT_7, TXTMCNT2296_4, SPAREO9, 
        CMDSMNXT_12, CMDSMNXT_3, SL_ET_ERR2723, TXDLCNT2426_1, SL_SP_ET_0, 
        TXDLCNT2418_6, CMDSTATE_13, NXTISTX, SPAREO0, SL_SP_E2648, 
        TXTMCNT2304_7, TXDLCNT_3, TXTMCNT2304_0, SL_SP_SC, TXDLCNT_4, 
        W4SOFGEN401, CMDSTATE_11, CMDSMNXT_4, SPAREO7, SL_SP_ET2642_1, 
        TEST_PACKET_T, SL_ACK_ERR2906, NXTISIDL, NEWCMD2004, TXDLCNT2418_1, 
        NXTISRCV, TXDLCNT2426_6, W4REPLY2010, SL_RXSPLIT, TXTMCNT2296_3, 
        ASKREPLY_3T, TXTMCNT_0, SPAREO5, CMDSTATE_10, CMDSTATE_6, 
        PHASENXT_CMD_SOF, n2356, TXDLCNT_6, ASKREPLY_2T, TXTMCNT2304_2, 
        TXTMCNT_2, TXTMCNT2296_1, CMDSMNXT_6, TXDLCNT2426_4, TX_PERIOD_P, 
        TXDLCNT2418_3, TXDLCNT2418_4, SL_SP_S2654, TXDLCNT2426_3, 
        TXTMCNT2296_6, TXSTART_D, PHASENXT_TERM, TXTMCNT_5, CMDSMNXT_8, 
        TXDLCNT_1, TX_PERIOD_P2529, TXTMCNT2304_5, TXDELAY, RCV_POWERUP_COND, 
        SPAREO2, TXTMCNT_4, TXTMCNT2296_7, TXTMOUT2366, TXDLCNT2426_2, 
        CMDSMNXT_9, TXDLCNT2418_5, SPAREO3, SL_SP_SC2660, SPAREO1_, 
        TXDELAY2488, TXDLCNT_0, ASKREPLY_PRE, PHASENXT_CMD_RXTOKEN, TXTMOUT, 
        ASKREPLY_T, TXTMCNT2304_4, RCV_POWERUP2134, TXDLCNT_7, TXTMCNT2304_3, 
        SPAREO4, CMDSTATE_0, CMDSMNXT_7, TXSTART_T, TXDLCNT2418_2, 
        TXDLCNT2426_5, TXTMCNT2296_0, TXTMCNT_3, n3260, n3263, n3264, n3265, 
        n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, 
        n3276, n3277, n3278, add_661_carry_6, add_661_carry_7, add_661_carry_2, 
        add_661_carry_5, add_661_carry_4, add_661_carry_3, n3300, n3301, n3302, 
        n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, 
        n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, 
        n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, 
        n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, 
        add_685_carry_6, add_685_carry_7, add_685_carry_2, add_685_carry_5, 
        add_685_carry_4, add_685_carry_3, n3342, n3343, n3344, n3345, n3346, 
        n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, 
        n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, 
        n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, 
        n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, 
        n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, 
        n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, 
        n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, 
        n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, 
        n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, 
        n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
        n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, 
        n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
        n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, 
        n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
        n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, 
        n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, 
        n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, 
        n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, 
        n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, 
        n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, 
        n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, 
        n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, 
        n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, 
        n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
        n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, 
        n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
        n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3615;
    zaoi211b SPARE632 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE635 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zoai21b SPARE634 ( .A(SPAREO0), .B(SPAREO8), .C(RCV_POWERUP_COND), .Y(
        SPAREO9) );
    zaoi211b SPARE633 ( .A(SPAREO4), .B(CURISTX), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zdffrb SPARE631 ( .CK(CLK60M), .D(SPAREO7), .R(TRST_), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE638 ( .A(SPAREO5), .Y(SPAREO6) );
    znr3b SPARE636 ( .A(SPAREO2), .B(NXTISTX), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE637 ( .A(SPAREO4), .Y(SPAREO5) );
    zdffrb SPARE630 ( .CK(CLK60M), .D(1'b0), .R(TRST_), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE639 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    znd2b U1083 ( .A(TXTMCNT_1), .B(n3334), .Y(n3307) );
    znr2b U1084 ( .A(TXTMCNT_0), .B(n3319), .Y(n3314) );
    zivb U1085 ( .A(TMOUT_PARM[0]), .Y(n3319) );
    znr2b U1086 ( .A(TXTMCNT_2), .B(n3336), .Y(n3337) );
    zivb U1087 ( .A(TMOUT_PARM[2]), .Y(n3336) );
    znr2b U1088 ( .A(TXTMCNT_1), .B(n3334), .Y(n3335) );
    zivb U1089 ( .A(TMOUT_PARM[1]), .Y(n3334) );
    znd2b U1090 ( .A(TXDLCNT_1), .B(n3376), .Y(n3349) );
    znr2b U1091 ( .A(TXDLCNT_0), .B(n3361), .Y(n3356) );
    zivb U1092 ( .A(TXDELAY_PARM[0]), .Y(n3361) );
    znr2b U1093 ( .A(TXDLCNT_2), .B(n3378), .Y(n3379) );
    zivb U1094 ( .A(TXDELAY_PARM[2]), .Y(n3378) );
    znr2b U1095 ( .A(TXDLCNT_1), .B(n3376), .Y(n3377) );
    zivb U1096 ( .A(TXDELAY_PARM[1]), .Y(n3376) );
    znd2b U1097 ( .A(n3313), .B(n3306), .Y(n3305) );
    znr2b U1098 ( .A(n3335), .B(n3337), .Y(n3313) );
    znd2b U1099 ( .A(n3314), .B(n3307), .Y(n3306) );
    znr2b U1100 ( .A(n3339), .B(n3333), .Y(n3312) );
    znr2b U1101 ( .A(TMOUT_PARM[2]), .B(n3338), .Y(n3339) );
    znr2b U1102 ( .A(TMOUT_PARM[3]), .B(n3332), .Y(n3333) );
    znr2b U1103 ( .A(TXTMCNT_4), .B(n3328), .Y(n3329) );
    zivb U1104 ( .A(TMOUT_PARM[4]), .Y(n3328) );
    znr2b U1105 ( .A(TXTMCNT_3), .B(n3326), .Y(n3327) );
    zivb U1106 ( .A(TMOUT_PARM[3]), .Y(n3326) );
    znd2b U1107 ( .A(n3355), .B(n3348), .Y(n3347) );
    znr2b U1108 ( .A(n3377), .B(n3379), .Y(n3355) );
    znd2b U1109 ( .A(n3356), .B(n3349), .Y(n3348) );
    znr2b U1110 ( .A(n3381), .B(n3375), .Y(n3354) );
    znr2b U1111 ( .A(TXDELAY_PARM[2]), .B(n3380), .Y(n3381) );
    znr2b U1112 ( .A(TXDELAY_PARM[3]), .B(n3374), .Y(n3375) );
    znr2b U1113 ( .A(TXDLCNT_4), .B(n3370), .Y(n3371) );
    zivb U1114 ( .A(TXDELAY_PARM[4]), .Y(n3370) );
    znr2b U1115 ( .A(TXDLCNT_3), .B(n3368), .Y(n3369) );
    zivb U1116 ( .A(TXDELAY_PARM[3]), .Y(n3368) );
    znd2b U1117 ( .A(n3311), .B(n3304), .Y(n3303) );
    znr2b U1118 ( .A(n3327), .B(n3329), .Y(n3311) );
    znd2b U1119 ( .A(n3312), .B(n3305), .Y(n3304) );
    znr2b U1120 ( .A(n3331), .B(n3325), .Y(n3310) );
    znr2b U1121 ( .A(TMOUT_PARM[4]), .B(n3330), .Y(n3331) );
    znr2b U1122 ( .A(TMOUT_PARM[5]), .B(n3324), .Y(n3325) );
    znr2b U1123 ( .A(TXTMCNT_5), .B(n3322), .Y(n3323) );
    zivb U1124 ( .A(TMOUT_PARM[5]), .Y(n3322) );
    znr2b U1125 ( .A(TXTMCNT_6), .B(n3320), .Y(n3321) );
    znd2b U1126 ( .A(n3353), .B(n3346), .Y(n3345) );
    znr2b U1127 ( .A(n3369), .B(n3371), .Y(n3353) );
    znd2b U1128 ( .A(n3354), .B(n3347), .Y(n3346) );
    znr2b U1129 ( .A(n3373), .B(n3367), .Y(n3352) );
    znr2b U1130 ( .A(TXDELAY_PARM[4]), .B(n3372), .Y(n3373) );
    znr2b U1131 ( .A(TXDELAY_PARM[5]), .B(n3366), .Y(n3367) );
    znr2b U1132 ( .A(TXDLCNT_5), .B(n3364), .Y(n3365) );
    zivb U1133 ( .A(TXDELAY_PARM[5]), .Y(n3364) );
    znr2b U1134 ( .A(TXDLCNT_6), .B(n3362), .Y(n3363) );
    zor2b U1135 ( .A(RXSETUP), .B(RXOUT), .Y(n3590) );
    zan2b U1136 ( .A(RXIN), .B(n3615), .Y(n3518) );
    znd2b U1137 ( .A(TXTMCNT_6), .B(n3320), .Y(n3316) );
    zivb U1138 ( .A(TMOUT_PARM[6]), .Y(n3320) );
    znd2b U1139 ( .A(n3309), .B(n3302), .Y(n3317) );
    znr2b U1140 ( .A(n3321), .B(n3323), .Y(n3309) );
    znd2b U1141 ( .A(n3310), .B(n3303), .Y(n3302) );
    znd2b U1142 ( .A(TXDLCNT_6), .B(n3362), .Y(n3358) );
    zivb U1143 ( .A(TXDELAY_PARM[6]), .Y(n3362) );
    znd2b U1144 ( .A(n3351), .B(n3344), .Y(n3359) );
    znr2b U1145 ( .A(n3363), .B(n3365), .Y(n3351) );
    znd2b U1146 ( .A(n3352), .B(n3345), .Y(n3344) );
    zao32b U1147 ( .A(n3571), .B(n3440), .C(n3499), .D(n3437), .E(n3391), .Y(
        n3484) );
    zivb U1148 ( .A(TD_PING), .Y(n3571) );
    zor2b U1149 ( .A(CMDSTATE_10), .B(n3453), .Y(n3530) );
    zoa22b U1150 ( .A(n3600), .B(n3555), .C(n3601), .D(n3545), .Y(n3599) );
    zmux21lb U1151 ( .A(n3518), .B(n3590), .S(SL_SP_SC), .Y(n3589) );
    zan2b U1152 ( .A(n3516), .B(n3517), .Y(n3419) );
    znd2b U1153 ( .A(n3300), .B(n3308), .Y(n3340) );
    znd2b U1154 ( .A(n3301), .B(n3315), .Y(n3300) );
    zivb U1155 ( .A(TMOUT_PARM[7]), .Y(n3308) );
    znd2b U1156 ( .A(TXTMCNT_7), .B(n3318), .Y(n3341) );
    znd2b U1157 ( .A(n3317), .B(n3316), .Y(n3318) );
    zivb U1158 ( .A(n3318), .Y(n3301) );
    zor2b U1159 ( .A(TXACK), .B(TXPING), .Y(n3529) );
    zivb U1160 ( .A(n3529), .Y(n3600) );
    zxo2b U1161 ( .A(n3442), .B(n3588), .Y(n3513) );
    zmux21lb U1162 ( .A(ASYNC_CMD[23]), .B(PERIOD_CMD[23]), .S(SL_PERIOD), .Y(
        n3588) );
    zxo2b U1163 ( .A(n3576), .B(n3597), .Y(n3512) );
    zmux21lb U1164 ( .A(ASYNC_CMD[22]), .B(PERIOD_CMD[22]), .S(SL_PERIOD), .Y(
        n3597) );
    zor2b U1165 ( .A(n3440), .B(n3538), .Y(n3496) );
    zivb U1166 ( .A(SP_SC), .Y(n3538) );
    zan2b U1167 ( .A(n3465), .B(n3466), .Y(n3464) );
    zivb U1168 ( .A(n3519), .Y(SL_PID[2]) );
    zor2b U1169 ( .A(RXSOF), .B(RXSPLIT), .Y(n3481) );
    zor2b U1170 ( .A(n3559), .B(n3557), .Y(n3558) );
    zivb U1171 ( .A(n3520), .Y(SL_PID[1]) );
    zivb U1172 ( .A(n3521), .Y(SL_PID[0]) );
    zor2b U1173 ( .A(n3516), .B(ISO), .Y(n3557) );
    zivb U1174 ( .A(n3557), .Y(n3492) );
    zan3b U1175 ( .A(TXTMOUT_EN), .B(n3501), .C(n3476), .Y(n3425) );
    zivb U1176 ( .A(NORMPKT), .Y(n3476) );
    zor2b U1177 ( .A(n3403), .B(n3556), .Y(n3493) );
    zor2b U1178 ( .A(n3566), .B(n3567), .Y(n3497) );
    zao21b U1179 ( .A(EOF1), .B(n3395), .C(n3270), .Y(n3415) );
    znd2b U1180 ( .A(n3611), .B(n3612), .Y(n3428) );
    zivb U1181 ( .A(n3593), .Y(n3559) );
    zor2b U1182 ( .A(NXTISRCV), .B(n3403), .Y(n3504) );
    zor2b U1183 ( .A(SP_SC), .B(n3440), .Y(n3535) );
    zivb U1184 ( .A(n3535), .Y(n3466) );
    zivb U1185 ( .A(RXSPLIT), .Y(n3573) );
    zan3b U1186 ( .A(n3507), .B(n3508), .C(n3509), .Y(n3506) );
    zivb U1187 ( .A(RXIN), .Y(n3507) );
    zxo2b U1188 ( .A(n3441), .B(SL_SP_E), .Y(n3511) );
    zxo2b U1189 ( .A(SL_SP_S), .B(n3587), .Y(n3510) );
    zmux21lb U1190 ( .A(n3595), .B(n3596), .S(RXIN), .Y(n3587) );
    znd2b U1191 ( .A(n3342), .B(n3350), .Y(n3382) );
    znd2b U1192 ( .A(n3343), .B(n3357), .Y(n3342) );
    zivb U1193 ( .A(TXDELAY_PARM[7]), .Y(n3350) );
    znd2b U1194 ( .A(TXDLCNT_7), .B(n3360), .Y(n3383) );
    znd2b U1195 ( .A(n3359), .B(n3358), .Y(n3360) );
    zivb U1196 ( .A(n3360), .Y(n3343) );
    zor2b U1197 ( .A(n3452), .B(n3453), .Y(CURISTX) );
    zor2b U1198 ( .A(TXSPLIT), .B(n3529), .Y(n3453) );
    zivb U1199 ( .A(n3453), .Y(n3601) );
    znr6b U1200 ( .A(n3275), .B(n3263), .C(n3264), .D(n3276), .E(n3481), .F(
        n3482), .Y(n3480) );
    zan3b U1201 ( .A(n3411), .B(n3487), .C(n3488), .Y(n3486) );
    zoai2x4b U1202 ( .A(n3606), .B(n3502), .C(n3607), .D(n3608), .E(n3609), 
        .F(n3543), .G(n3554), .H(n3556), .Y(n3605) );
    zivb U1203 ( .A(n3517), .Y(n3607) );
    zor2b U1204 ( .A(TXOUT), .B(TXSETUP), .Y(n3517) );
    zivb U1205 ( .A(n3524), .Y(n3608) );
    zor2b U1206 ( .A(TXSOF), .B(TXIN), .Y(n3524) );
    zivb U1207 ( .A(n3525), .Y(n3609) );
    zor2b U1208 ( .A(n3524), .B(n3517), .Y(n3525) );
    zivb U1209 ( .A(EOF1), .Y(n3556) );
    zivb U1210 ( .A(n3554), .Y(n3499) );
    zao32b U1211 ( .A(n3270), .B(n3423), .C(PKRVEND), .D(n3271), .E(PKTXEND), 
        .Y(n3569) );
    zivb U1212 ( .A(n3569), .Y(n3611) );
    zmux21lb U1213 ( .A(n3591), .B(EOF2), .S(EOF1), .Y(n3485) );
    zoa211b U1214 ( .A(TXDELAY_EN), .B(n3475), .C(n3592), .D(n3593), .Y(n3591)
         );
    zor2b U1215 ( .A(n3539), .B(n3418), .Y(n3495) );
    zivc U1216 ( .A(n3577), .Y(n3563) );
    zor2b U1217 ( .A(CMDSTATE_13), .B(CMDSTATE_11), .Y(n3522) );
    zor2b U1218 ( .A(CMDSTATE_14), .B(n3530), .Y(n3531) );
    zan2b U1219 ( .A(n3478), .B(n3479), .Y(n3477) );
    zor2b U1220 ( .A(CMDSTATE_5), .B(n3525), .Y(n3452) );
    zor2b U1221 ( .A(CMDSTATE_0), .B(n3445), .Y(n3523) );
    zan3b U1222 ( .A(n3472), .B(n3473), .C(n3474), .Y(n3471) );
    zoa22b U1223 ( .A(n3552), .B(n3467), .C(n3528), .D(n3560), .Y(n3472) );
    zoa211b U1224 ( .A(n3602), .B(n3468), .C(n3599), .D(n3603), .Y(n3473) );
    zivb U1225 ( .A(n3530), .Y(n3602) );
    zxo2b U1226 ( .A(n3580), .B(n3581), .Y(n3474) );
    zivb U1227 ( .A(n3522), .Y(n3580) );
    zivb U1228 ( .A(n3531), .Y(n3581) );
    zivb U1229 ( .A(n3463), .Y(n3449) );
    zivb U1230 ( .A(n3462), .Y(n3450) );
    zivb U1231 ( .A(n3461), .Y(n3456) );
    zxo2b U1232 ( .A(RXPID[0]), .B(SL_MAXLEN[8]), .Y(n3583) );
    zxo2b U1233 ( .A(RXPID[2]), .B(SL_MAXLEN[10]), .Y(n3582) );
    zxo2b U1234 ( .A(RXPID[3]), .B(n3586), .Y(n3585) );
    zivb U1235 ( .A(n3596), .Y(n3586) );
    zmux21lb U1236 ( .A(ASYNC_CMD[19]), .B(PERIOD_CMD[19]), .S(SL_PERIOD), .Y(
        n3596) );
    zxo2b U1237 ( .A(RXPID[1]), .B(SL_MAXLEN[9]), .Y(n3584) );
    zor2b U1238 ( .A(n3542), .B(n3545), .Y(n3572) );
    zan2b U1239 ( .A(n3265), .B(TXTMCNT2296_7), .Y(TXTMCNT2304_7) );
    zxo2b U1240 ( .A(add_661_carry_7), .B(TXTMCNT_7), .Y(TXTMCNT2296_7) );
    zan2b U1241 ( .A(TXTMCNT2296_6), .B(n3265), .Y(TXTMCNT2304_6) );
    zhadrb add_661_U1_1_6 ( .A(TXTMCNT_6), .B(add_661_carry_6), .CO(
        add_661_carry_7), .S(TXTMCNT2296_6) );
    zan2b U1242 ( .A(TXTMCNT2296_5), .B(n3265), .Y(TXTMCNT2304_5) );
    zhadrb add_661_U1_1_5 ( .A(TXTMCNT_5), .B(add_661_carry_5), .CO(
        add_661_carry_6), .S(TXTMCNT2296_5) );
    zan2b U1243 ( .A(TXTMCNT2296_4), .B(n3265), .Y(TXTMCNT2304_4) );
    zhadrb add_661_U1_1_4 ( .A(TXTMCNT_4), .B(add_661_carry_4), .CO(
        add_661_carry_5), .S(TXTMCNT2296_4) );
    zan2b U1244 ( .A(TXTMCNT2296_3), .B(n3265), .Y(TXTMCNT2304_3) );
    zhadrb add_661_U1_1_3 ( .A(TXTMCNT_3), .B(add_661_carry_3), .CO(
        add_661_carry_4), .S(TXTMCNT2296_3) );
    zan2b U1245 ( .A(TXTMCNT2296_2), .B(n3265), .Y(TXTMCNT2304_2) );
    zhadrb add_661_U1_1_2 ( .A(TXTMCNT_2), .B(add_661_carry_2), .CO(
        add_661_carry_3), .S(TXTMCNT2296_2) );
    zan2b U1246 ( .A(TXTMCNT2296_1), .B(n3265), .Y(TXTMCNT2304_1) );
    zhadrb add_661_U1_1_1 ( .A(TXTMCNT_1), .B(TXTMCNT_0), .CO(add_661_carry_2), 
        .S(TXTMCNT2296_1) );
    zan2b U1247 ( .A(TXTMCNT2296_0), .B(n3265), .Y(TXTMCNT2304_0) );
    zan2b U1248 ( .A(n3266), .B(TXDLCNT2418_7), .Y(TXDLCNT2426_7) );
    zxo2b U1249 ( .A(add_685_carry_7), .B(TXDLCNT_7), .Y(TXDLCNT2418_7) );
    zan2b U1250 ( .A(TXDLCNT2418_6), .B(n3266), .Y(TXDLCNT2426_6) );
    zhadrb add_685_U1_1_6 ( .A(TXDLCNT_6), .B(add_685_carry_6), .CO(
        add_685_carry_7), .S(TXDLCNT2418_6) );
    zan2b U1251 ( .A(TXDLCNT2418_5), .B(n3266), .Y(TXDLCNT2426_5) );
    zhadrb add_685_U1_1_5 ( .A(TXDLCNT_5), .B(add_685_carry_5), .CO(
        add_685_carry_6), .S(TXDLCNT2418_5) );
    zan2b U1252 ( .A(TXDLCNT2418_4), .B(n3266), .Y(TXDLCNT2426_4) );
    zhadrb add_685_U1_1_4 ( .A(TXDLCNT_4), .B(add_685_carry_4), .CO(
        add_685_carry_5), .S(TXDLCNT2418_4) );
    zan2b U1253 ( .A(TXDLCNT2418_3), .B(n3266), .Y(TXDLCNT2426_3) );
    zhadrb add_685_U1_1_3 ( .A(TXDLCNT_3), .B(add_685_carry_3), .CO(
        add_685_carry_4), .S(TXDLCNT2418_3) );
    zan2b U1254 ( .A(TXDLCNT2418_2), .B(n3266), .Y(TXDLCNT2426_2) );
    zhadrb add_685_U1_1_2 ( .A(TXDLCNT_2), .B(add_685_carry_2), .CO(
        add_685_carry_3), .S(TXDLCNT2418_2) );
    zan2b U1255 ( .A(TXDLCNT2418_1), .B(n3266), .Y(TXDLCNT2426_1) );
    zhadrb add_685_U1_1_1 ( .A(TXDLCNT_1), .B(TXDLCNT_0), .CO(add_685_carry_2), 
        .S(TXDLCNT2418_1) );
    zan2b U1256 ( .A(TXDLCNT2418_0), .B(n3266), .Y(TXDLCNT2426_0) );
    zao22b U1257 ( .A(SL_SP_ET_1), .B(n3267), .C(RXADDRF[18]), .D(n3272), .Y(
        SL_SP_ET2642_1) );
    zao22b U1258 ( .A(SL_SP_ET_0), .B(n3267), .C(RXADDRF[17]), .D(n3272), .Y(
        SL_SP_ET2642_0) );
    zivb U1259 ( .A(TD_IN), .Y(n3410) );
    zivb U1260 ( .A(CMDSMNXT_2), .Y(n3433) );
    zivb U1261 ( .A(n3568), .Y(n3501) );
    zivb U1262 ( .A(CMDSMNXT_12), .Y(n3434) );
    zao32b U1263 ( .A(TEST_PACKET), .B(n3411), .C(MAC_CMDSTART), .D(n3264), 
        .E(n3394), .Y(n3384) );
    zan3b U1264 ( .A(n3496), .B(n3497), .C(n3391), .Y(n3385) );
    zivb U1265 ( .A(CMDSMNXT_5), .Y(n3436) );
    zao21b U1266 ( .A(EOFTERM), .B(n3455), .C(PHASENXT_TERM), .Y(EOFTERM2247)
         );
    zivb U1267 ( .A(SOFGEN), .Y(n3455) );
    zao32b U1268 ( .A(n3430), .B(MAC_EOT), .C(n3447), .D(n3260), .E(
        MAC_SLAVE_ACT), .Y(NEWCMD2004) );
    zao21b U1269 ( .A(TX_PERIOD_P), .B(n3403), .C(TXSTART), .Y(TX_PERIOD_P2529
        ) );
    zivb U1270 ( .A(TD_SETUP), .Y(n3389) );
    zivb U1271 ( .A(CMDSMNXT_4), .Y(n3435) );
    zivb U1272 ( .A(n3387), .Y(n3566) );
    zao22b U1273 ( .A(SL_SP_E), .B(n3267), .C(RXADDRF[16]), .D(n3272), .Y(
        SL_SP_E2648) );
    zor2b U1274 ( .A(CMDSTATE_6), .B(DATAIN), .Y(n3445) );
    zivb U1275 ( .A(n3445), .Y(n3606) );
    zan2b U1276 ( .A(PKTXEND), .B(NXTISRCV), .Y(W4REPLY2010) );
    zor2b U1277 ( .A(EOF1), .B(n3498), .Y(n3388) );
    zivb U1278 ( .A(TD_OUT), .Y(n3439) );
    zivb U1279 ( .A(CMDSMNXT_3), .Y(n3432) );
    zivb U1280 ( .A(n3438), .Y(n3567) );
    znd2b U1281 ( .A(n3341), .B(n3340), .Y(n2356) );
    zao22b U1282 ( .A(n3437), .B(n3403), .C(n3274), .D(TD_SPLIT), .Y(
        CMDSMNXT_8) );
    zivb U1283 ( .A(n3500), .Y(n3437) );
    zivb U1284 ( .A(CMDSMNXT_8), .Y(n3429) );
    zao22b U1285 ( .A(n3267), .B(SL_SP_SC), .C(RXADDRF[7]), .D(n3272), .Y(
        SL_SP_SC2660) );
    zao22b U1286 ( .A(SL_SP_S), .B(n3267), .C(RXADDRF[15]), .D(n3272), .Y(
        SL_SP_S2654) );
    zivb U1287 ( .A(n3574), .Y(n3575) );
    zao32b U1288 ( .A(n3411), .B(n3412), .C(n3413), .D(n3414), .E(n3403), .Y(
        PHASENXT_CMD_SOF) );
    zor2b U1289 ( .A(SOFGEN), .B(W4SOFGEN), .Y(n3412) );
    zoai21b U1290 ( .A(MAC_SLAVE_ACT), .B(TEST_PACKET), .C(MAC_CMDSTART), .Y(
        n3413) );
    zivb U1291 ( .A(n3565), .Y(n3414) );
    zivb U1292 ( .A(PHASENXT_CMD_SOF), .Y(n3430) );
    zivb U1293 ( .A(n3412), .Y(n3488) );
    zor2b U1294 ( .A(n3448), .B(SL_ET_ERR), .Y(SL_ET_ERR2723) );
    zivb U1295 ( .A(n3496), .Y(n3516) );
    zivb U1296 ( .A(n3494), .Y(n3393) );
    zivf U1297 ( .A(n3418), .Y(n3544) );
    zor2b U1298 ( .A(SL_ACK_ERR), .B(n3451), .Y(SL_ACK_ERR2906) );
    zmux21lb U1299 ( .A(n3598), .B(n3572), .S(RXACK), .Y(n3451) );
    zao21b U1300 ( .A(W4SOFGEN), .B(CMDSTATE_0), .C(SOFGEN), .Y(W4SOFGEN401)
         );
    znr8b U1301 ( .A(n3446), .B(CMDSMNXT_14), .C(PHASENXT_TERM), .D(
        CMDSMNXT_13), .E(NXTISIDL), .F(n3260), .G(TXSTART), .H(
        PHASENXT_CMD_RXTOKEN), .Y(TXSTART_D) );
    zao32b U1302 ( .A(n3426), .B(n3427), .C(n3423), .D(TXDELAY_EN), .E(n3428), 
        .Y(CMDSMNXT_14) );
    zivb U1303 ( .A(n3561), .Y(n3426) );
    zivb U1304 ( .A(EOF2), .Y(n3423) );
    zao32b U1305 ( .A(PKRVEND), .B(EOF2), .C(n3415), .D(n3416), .E(n3417), .Y(
        PHASENXT_TERM) );
    zivb U1306 ( .A(n3493), .Y(n3416) );
    zao32b U1307 ( .A(n3421), .B(n3422), .C(n3423), .D(n3424), .E(n3425), .Y(
        CMDSMNXT_13) );
    zivb U1308 ( .A(n3562), .Y(n3421) );
    zivb U1309 ( .A(n3558), .Y(n3424) );
    zivb U1310 ( .A(n3481), .Y(n3579) );
    zor2b U1311 ( .A(n3454), .B(SL_DATA_PIDERR), .Y(SL_DATA_PIDERR2868) );
    zan3b U1312 ( .A(PKRVEND), .B(DATAIN), .C(n3514), .Y(n3454) );
    zivb U1313 ( .A(n3482), .Y(n3394) );
    zor2b U1314 ( .A(n3546), .B(n3390), .Y(n3482) );
    zivb U1315 ( .A(RXOUT), .Y(n3509) );
    zivb U1316 ( .A(RXSETUP), .Y(n3508) );
    zan2b U1317 ( .A(n3465), .B(n3535), .Y(n3396) );
    zivb U1318 ( .A(n3409), .Y(n3465) );
    zivb U1319 ( .A(n3539), .Y(n3391) );
    zor2b U1320 ( .A(EOF1), .B(n3403), .Y(n3539) );
    zao21b U1321 ( .A(SL_RXSPLIT), .B(n3459), .C(n3272), .Y(SL_RXSPLIT2598) );
    zor2b U1322 ( .A(n3458), .B(SL_SE_ERR), .Y(SL_SE_ERR2808) );
    zao32b U1323 ( .A(TD_PING), .B(n3440), .C(n3274), .D(n3268), .E(n3403), 
        .Y(CMDSMNXT_9) );
    zivb U1324 ( .A(TD_SPLIT), .Y(n3440) );
    zivb U1325 ( .A(MAC_CMDSTART), .Y(n3487) );
    zivb U1326 ( .A(CMDSMNXT_9), .Y(n3431) );
    znd2b U1327 ( .A(n3383), .B(n3382), .Y(n2478) );
    zivb U1328 ( .A(n3546), .Y(n3406) );
    zivb U1329 ( .A(PKRVEND), .Y(n3390) );
    zivb U1330 ( .A(n3551), .Y(n3469) );
    zivb U1331 ( .A(n3553), .Y(n3411) );
    zivb U1332 ( .A(TEST_PACKET), .Y(n3470) );
    zmux21lb U1333 ( .A(n3594), .B(n3471), .S(n3477), .Y(n3397) );
    zivb U1334 ( .A(n3532), .Y(n3594) );
    zoai2x4b U1335 ( .A(n3561), .B(n3427), .C(n3479), .D(n3478), .E(n3562), 
        .F(n3422), .G(n3403), .H(n3565), .Y(n3399) );
    zivb U1336 ( .A(n3523), .Y(n3479) );
    zivb U1337 ( .A(n3452), .Y(n3478) );
    zivb U1338 ( .A(PKTXEND), .Y(n3403) );
    zan2b U1339 ( .A(n3490), .B(n3269), .Y(n3400) );
    zivb U1340 ( .A(n3495), .Y(n3490) );
    zan3b U1341 ( .A(n3395), .B(PKRVEND), .C(n3485), .Y(n3401) );
    zivb U1342 ( .A(n3550), .Y(n3395) );
    zivb U1343 ( .A(TXDELAY_EN), .Y(n3570) );
    zivb U1344 ( .A(NXTISIDL), .Y(n3447) );
    zivb U1345 ( .A(n3514), .Y(SL_TOGMATCH) );
    zivb U1346 ( .A(n3459), .Y(MAC_EOT) );
    zor2b U1347 ( .A(W4SOFGEN), .B(n3502), .Y(n3459) );
    zivb U1348 ( .A(n3572), .Y(RXTOKENPHASE) );
    zan2b U1349 ( .A(DATM), .B(CMDSTATE_5), .Y(TXMDATA) );
    zan2b U1350 ( .A(DAT2), .B(CMDSTATE_5), .Y(TXDATA2) );
    zan2b U1351 ( .A(DAT1), .B(CMDSTATE_5), .Y(TXDATA1) );
    zor2b U1352 ( .A(n3457), .B(SL_TXDATASEL[2]), .Y(TXDATA0) );
    zivb U1353 ( .A(MAC_SLAVE_ACT), .Y(n3542) );
    zdffqrb TXTMCNT_reg_7 ( .CK(CLK60M), .D(TXTMCNT2304_7), .R(TRST_), .Q(
        TXTMCNT_7) );
    zivb U1354 ( .A(TXTMCNT_7), .Y(n3315) );
    zdffqrb TXTMCNT_reg_6 ( .CK(CLK60M), .D(TXTMCNT2304_6), .R(TRST_), .Q(
        TXTMCNT_6) );
    zdffqrb TXTMCNT_reg_5 ( .CK(CLK60M), .D(TXTMCNT2304_5), .R(TRST_), .Q(
        TXTMCNT_5) );
    zivb U1355 ( .A(TXTMCNT_5), .Y(n3324) );
    zdffqrb TXTMCNT_reg_4 ( .CK(CLK60M), .D(TXTMCNT2304_4), .R(TRST_), .Q(
        TXTMCNT_4) );
    zivb U1356 ( .A(TXTMCNT_4), .Y(n3330) );
    zdffqrb TXTMCNT_reg_3 ( .CK(CLK60M), .D(TXTMCNT2304_3), .R(TRST_), .Q(
        TXTMCNT_3) );
    zivb U1357 ( .A(TXTMCNT_3), .Y(n3332) );
    zdffqrb TXTMCNT_reg_2 ( .CK(CLK60M), .D(TXTMCNT2304_2), .R(TRST_), .Q(
        TXTMCNT_2) );
    zivb U1358 ( .A(TXTMCNT_2), .Y(n3338) );
    zdffqrb TXTMCNT_reg_1 ( .CK(CLK60M), .D(TXTMCNT2304_1), .R(TRST_), .Q(
        TXTMCNT_1) );
    zdffqrb TXTMCNT_reg_0 ( .CK(CLK60M), .D(TXTMCNT2304_0), .R(TRST_), .Q(
        TXTMCNT_0) );
    zivb U1359 ( .A(TXTMCNT_0), .Y(TXTMCNT2296_0) );
    zdffqrb TXDLCNT_reg_7 ( .CK(CLK60M), .D(TXDLCNT2426_7), .R(TRST_), .Q(
        TXDLCNT_7) );
    zivb U1360 ( .A(TXDLCNT_7), .Y(n3357) );
    zdffqrb TXDLCNT_reg_6 ( .CK(CLK60M), .D(TXDLCNT2426_6), .R(TRST_), .Q(
        TXDLCNT_6) );
    zdffqrb TXDLCNT_reg_5 ( .CK(CLK60M), .D(TXDLCNT2426_5), .R(TRST_), .Q(
        TXDLCNT_5) );
    zivb U1361 ( .A(TXDLCNT_5), .Y(n3366) );
    zdffqrb TXDLCNT_reg_4 ( .CK(CLK60M), .D(TXDLCNT2426_4), .R(TRST_), .Q(
        TXDLCNT_4) );
    zivb U1362 ( .A(TXDLCNT_4), .Y(n3372) );
    zdffqrb TXDLCNT_reg_3 ( .CK(CLK60M), .D(TXDLCNT2426_3), .R(TRST_), .Q(
        TXDLCNT_3) );
    zivb U1363 ( .A(TXDLCNT_3), .Y(n3374) );
    zdffqrb TXDLCNT_reg_2 ( .CK(CLK60M), .D(TXDLCNT2426_2), .R(TRST_), .Q(
        TXDLCNT_2) );
    zivb U1364 ( .A(TXDLCNT_2), .Y(n3380) );
    zdffqrb TXDLCNT_reg_1 ( .CK(CLK60M), .D(TXDLCNT2426_1), .R(TRST_), .Q(
        TXDLCNT_1) );
    zdffqrb TXDLCNT_reg_0 ( .CK(CLK60M), .D(TXDLCNT2426_0), .R(TRST_), .Q(
        TXDLCNT_0) );
    zivb U1365 ( .A(TXDLCNT_0), .Y(TXDLCNT2418_0) );
    zdffqrb_ SL_SP_ET_reg_1 ( .CK(CLK60M), .D(SL_SP_ET2642_1), .R(TRST_), .Q(
        SL_SP_ET_1) );
    zivb U1366 ( .A(SL_SP_ET_1), .Y(n3442) );
    zdffqrb_ SL_SP_ET_reg_0 ( .CK(CLK60M), .D(SL_SP_ET2642_0), .R(TRST_), .Q(
        SL_SP_ET_0) );
    zivb U1367 ( .A(SL_SP_ET_0), .Y(n3576) );
    zdffqrb_ CMDSTATE_reg_2 ( .CK(CLK60M), .D(CMDSMNXT_2), .R(TRST_), .Q(TXIN)
         );
    zivb U1368 ( .A(TXIN), .Y(n3534) );
    zdffqrb_ CMDSTATE_reg_12 ( .CK(CLK60M), .D(CMDSMNXT_12), .R(TRST_), .Q(
        TXACK) );
    zivb U1369 ( .A(TXACK), .Y(n3560) );
    zdffqrb_ CMDSTATE_reg_15 ( .CK(CLK60M), .D(PHASENXT_TERM), .R(TRST_), .Q(
        CMDSTATE_15) );
    zivb U1370 ( .A(CMDSTATE_15), .Y(n3603) );
    zdffqrb_ CMDSTATE_reg_5 ( .CK(CLK60M), .D(CMDSMNXT_5), .R(TRST_), .Q(
        CMDSTATE_5) );
    zivb U1371 ( .A(CMDSTATE_5), .Y(n3543) );
    zdffqrb TXSTART_reg ( .CK(CLK60M), .D(TXSTART_T), .R(TRST_), .Q(TXSTART)
         );
    zdffqrb_ EOFTERM_reg ( .CK(CLK60M), .D(EOFTERM2247), .R(TRST_), .Q(EOFTERM
        ) );
    zdffqrb_ NEWCMD_reg ( .CK(CLK60M), .D(NEWCMD2004), .R(TRST_), .Q(NEWCMD)
         );
    zdffqrb_ TX_PERIOD_P_reg ( .CK(CLK60M), .D(TX_PERIOD_P2529), .R(TRST_), 
        .Q(TX_PERIOD_P) );
    zdffqrb_ CMDSTATE_reg_4 ( .CK(CLK60M), .D(CMDSMNXT_4), .R(TRST_), .Q(
        TXSETUP) );
    zivb U1372 ( .A(TXSETUP), .Y(n3536) );
    zdffqrb_ CMDSTATE_reg_14 ( .CK(CLK60M), .D(CMDSMNXT_14), .R(TRST_), .Q(
        CMDSTATE_14) );
    zivb U1373 ( .A(CMDSTATE_14), .Y(n3468) );
    zdffqrb_ SL_SP_E_reg ( .CK(CLK60M), .D(SL_SP_E2648), .R(TRST_), .Q(SL_SP_E
        ) );
    zdffqrb_ ASKREPLY_PRE_reg ( .CK(CLK60M), .D(NXTISRCV), .R(TRST_), .Q(
        ASKREPLY_PRE) );
    zdffqrb_ TEST_PACKET_T_reg ( .CK(CLK60M), .D(TEST_PACKET), .R(TRST_), .Q(
        TEST_PACKET_T) );
    zdffqrb_ RCV_POWERUP_reg ( .CK(CLK60M), .D(RCV_POWERUP2134), .R(TRST_), 
        .Q(RCV_POWERUP) );
    zdffqrb_ CMDSTATE_reg_13 ( .CK(CLK60M), .D(CMDSMNXT_13), .R(TRST_), .Q(
        CMDSTATE_13) );
    zivb U1374 ( .A(CMDSTATE_13), .Y(n3467) );
    zdffqrb_ W4REPLY_reg ( .CK(CLK60M), .D(W4REPLY2010), .R(TRST_), .Q(W4REPLY
        ) );
    zdffqrb_ CMDSTATE_reg_3 ( .CK(CLK60M), .D(CMDSMNXT_3), .R(TRST_), .Q(TXOUT
        ) );
    zivb U1375 ( .A(TXOUT), .Y(n3537) );
    zdffqrb TXTMOUT_reg ( .CK(CLK60M), .D(TXTMOUT2366), .R(TRST_), .Q(TXTMOUT)
         );
    zivb U1376 ( .A(TXTMOUT), .Y(n3422) );
    zdffqrb_ CMDSTATE_reg_8 ( .CK(CLK60M), .D(CMDSMNXT_8), .R(TRST_), .Q(
        TXSPLIT) );
    zivb U1377 ( .A(TXSPLIT), .Y(n3555) );
    zdffqrb_ SL_SP_SC_reg ( .CK(CLK60M), .D(SL_SP_SC2660), .R(TRST_), .Q(
        SL_SP_SC) );
    zivb U1378 ( .A(SL_SP_SC), .Y(n3547) );
    zdffqrb_ SL_SP_S_reg ( .CK(CLK60M), .D(SL_SP_S2654), .R(TRST_), .Q(SL_SP_S
        ) );
    zdffqrb_ CMDSTATE_reg_1 ( .CK(CLK60M), .D(PHASENXT_CMD_SOF), .R(TRST_), 
        .Q(TXSOF) );
    zivb U1379 ( .A(TXSOF), .Y(n3564) );
    zdffqrb_ SL_ET_ERR_reg ( .CK(CLK60M), .D(SL_ET_ERR2723), .R(TRST_), .Q(
        SL_ET_ERR) );
    zdffqrb_ CMDSTATE_reg_11 ( .CK(CLK60M), .D(n3260), .R(TRST_), .Q(
        CMDSTATE_11) );
    zivb U1380 ( .A(CMDSTATE_11), .Y(n3552) );
    zdffqrb_ CMDSTATE_reg_6 ( .CK(CLK60M), .D(CMDSMNXT_6), .R(TRST_), .Q(
        CMDSTATE_6) );
    zivb U1381 ( .A(CMDSTATE_6), .Y(n3541) );
    zdffqrb_ SL_ACK_ERR_reg ( .CK(CLK60M), .D(SL_ACK_ERR2906), .R(TRST_), .Q(
        SL_ACK_ERR) );
    zdffqrb W4SOFGEN_reg ( .CK(CLK60M), .D(W4SOFGEN401), .R(TRST_), .Q(
        W4SOFGEN) );
    zivb U1382 ( .A(W4SOFGEN), .Y(n3503) );
    zdffqrb_ TXSTART_T_reg ( .CK(CLK60M), .D(TXSTART_D), .R(TRST_), .Q(
        TXSTART_T) );
    zdffqrb_ SL_DATA_PIDERR_reg ( .CK(CLK60M), .D(SL_DATA_PIDERR2868), .R(
        TRST_), .Q(SL_DATA_PIDERR) );
    zdffqrb_ CMDSTATE_reg_7 ( .CK(CLK60M), .D(CMDSMNXT_7), .R(TRST_), .Q(
        DATAIN) );
    zivb U1383 ( .A(DATAIN), .Y(n3549) );
    zdffqrb_ ASKREPLY_2T_reg ( .CK(CLK60M), .D(ASKREPLY_T), .R(TRST_), .Q(
        ASKREPLY_2T) );
    zdffqrb_ SL_RXSPLIT_reg ( .CK(CLK60M), .D(SL_RXSPLIT2598), .R(TRST_), .Q(
        SL_RXSPLIT) );
    zivb U1384 ( .A(SL_RXSPLIT), .Y(n3548) );
    zdffqrb_ SL_SE_ERR_reg ( .CK(CLK60M), .D(SL_SE_ERR2808), .R(TRST_), .Q(
        SL_SE_ERR) );
    zdffrb_ CMDSTATE_reg_9 ( .CK(CLK60M), .D(CMDSMNXT_9), .R(TRST_), .Q(TXPING
        ), .QN(n3528) );
    zdffqrb TXDELAY_reg ( .CK(CLK60M), .D(TXDELAY2488), .R(TRST_), .Q(TXDELAY)
         );
    zivb U1385 ( .A(TXDELAY), .Y(n3427) );
    zdffqrb_ ASKREPLY_3T_reg ( .CK(CLK60M), .D(ASKREPLY_2T), .R(TRST_), .Q(
        ASKREPLY_3T) );
    zdffqrb_ ASKREPLY_T_reg ( .CK(CLK60M), .D(ASKREPLY_PRE), .R(TRST_), .Q(
        ASKREPLY_T) );
    zdffqrb_ CMDSTATE_reg_10 ( .CK(CLK60M), .D(PHASENXT_CMD_RXTOKEN), .R(TRST_
        ), .Q(CMDSTATE_10) );
    zivb U1386 ( .A(CMDSTATE_10), .Y(n3545) );
    zdffqsb_ CMDSTATE_reg_0 ( .CK(CLK60M), .D(NXTISIDL), .S(TRST_), .Q(
        CMDSTATE_0) );
    zivb U1387 ( .A(CMDSTATE_0), .Y(n3502) );
    zivc U1388 ( .A(RXADDRF[0]), .Y(n3615) );
    znr2b U1389 ( .A(n3579), .B(n3482), .Y(n3260) );
    znr2b U1390 ( .A(n3542), .B(n3543), .Y(SL_TXDATASEL[2]) );
    zan2b U1391 ( .A(ASKREPLY_PRE), .B(ASKREPLY_3T), .Y(ASKREPLY) );
    znr3b U1392 ( .A(n3589), .B(n3548), .C(n3559), .Y(n3263) );
    zaoi211b U1393 ( .A(SL_RXSPLIT), .B(n3547), .C(n3507), .D(n3559), .Y(n3264
        ) );
    znr2b U1394 ( .A(TXTMOUT), .B(n3467), .Y(n3265) );
    znr2b U1395 ( .A(TXDELAY), .B(n3468), .Y(n3266) );
    znr2b U1396 ( .A(MAC_EOT), .B(n3575), .Y(n3267) );
    znr4b U1397 ( .A(TXACK), .B(TXSPLIT), .C(n3528), .D(n3527), .Y(n3268) );
    znr4b U1398 ( .A(n3523), .B(n3525), .C(n3543), .D(n3532), .Y(n3269) );
    znr3b U1399 ( .A(DATAIN), .B(n3541), .C(n3540), .Y(n3270) );
    znr4b U1400 ( .A(TXPING), .B(TXSPLIT), .C(n3560), .D(n3527), .Y(n3271) );
    znr2b U1401 ( .A(MAC_EOT), .B(n3574), .Y(n3272) );
    znr3b U1402 ( .A(n3463), .B(n3462), .C(n3461), .Y(n3273) );
    znr3b U1403 ( .A(EOF1), .B(n3487), .C(n3554), .Y(n3274) );
    zaoi22b U1404 ( .A(SL_RXSPLIT), .B(SL_SP_SC), .C(n3509), .D(n3508), .Y(
        n3275) );
    zan2b U1405 ( .A(RXPING), .B(n3593), .Y(n3276) );
    znr4b U1406 ( .A(n3506), .B(n3390), .C(n3548), .D(n3572), .Y(n3277) );
    znr2b U1407 ( .A(n3273), .B(n3542), .Y(n3278) );
    zmux21hb U1408 ( .A(ASYNC_CMD[27]), .B(PERIOD_CMD[27]), .S(SL_PERIOD), .Y(
        SL_PID[3]) );
    zmux21hb U1409 ( .A(ASYNC_CMD[20]), .B(PERIOD_CMD[20]), .S(n3613), .Y(
        SL_TXDATASEL[0]) );
    zmux21hb U1410 ( .A(ASYNC_CMD[18]), .B(PERIOD_CMD[18]), .S(SL_PERIOD), .Y(
        SL_MAXLEN[10]) );
    zmux21hb U1411 ( .A(ASYNC_CMD[16]), .B(PERIOD_CMD[16]), .S(n3613), .Y(
        SL_MAXLEN[8]) );
    zmux21hb U1412 ( .A(ASYNC_CMD[17]), .B(PERIOD_CMD[17]), .S(SL_PERIOD), .Y(
        SL_MAXLEN[9]) );
    zivc U1413 ( .A(n3615), .Y(n3613) );
    zivb U1414 ( .A(n3615), .Y(SL_PERIOD) );
    zbfb U1415 ( .A(SL_CRC16[0]), .Y(SL_TXFIXDATA[0]) );
    zmux21hb U1416 ( .A(ASYNC_CMD[0]), .B(PERIOD_CMD[0]), .S(n3613), .Y(
        SL_CRC16[0]) );
    zbfb U1417 ( .A(SL_CRC16[1]), .Y(SL_TXFIXDATA[1]) );
    zmux21hb U1418 ( .A(ASYNC_CMD[1]), .B(PERIOD_CMD[1]), .S(n3613), .Y(
        SL_CRC16[1]) );
    zbfb U1419 ( .A(SL_CRC16[2]), .Y(SL_TXFIXDATA[2]) );
    zmux21hb U1420 ( .A(ASYNC_CMD[2]), .B(PERIOD_CMD[2]), .S(n3613), .Y(
        SL_CRC16[2]) );
    zbfb U1421 ( .A(SL_CRC16[3]), .Y(SL_TXFIXDATA[3]) );
    zmux21hb U1422 ( .A(ASYNC_CMD[3]), .B(PERIOD_CMD[3]), .S(n3613), .Y(
        SL_CRC16[3]) );
    zbfb U1423 ( .A(SL_CRC16[4]), .Y(SL_TXFIXDATA[4]) );
    zmux21hb U1424 ( .A(ASYNC_CMD[4]), .B(PERIOD_CMD[4]), .S(n3613), .Y(
        SL_CRC16[4]) );
    zbfb U1425 ( .A(SL_CRC16[5]), .Y(SL_TXFIXDATA[5]) );
    zmux21hb U1426 ( .A(ASYNC_CMD[5]), .B(PERIOD_CMD[5]), .S(SL_PERIOD), .Y(
        SL_CRC16[5]) );
    zbfb U1427 ( .A(SL_CRC16[6]), .Y(SL_TXFIXDATA[6]) );
    zmux21hb U1428 ( .A(ASYNC_CMD[6]), .B(PERIOD_CMD[6]), .S(SL_PERIOD), .Y(
        SL_CRC16[6]) );
    zbfb U1429 ( .A(SL_CRC16[7]), .Y(SL_TXFIXDATA[7]) );
    zmux21hb U1430 ( .A(ASYNC_CMD[7]), .B(PERIOD_CMD[7]), .S(SL_PERIOD), .Y(
        SL_CRC16[7]) );
    zbfb U1431 ( .A(SL_CRC16[8]), .Y(SL_MAXLEN[0]) );
    zmux21hb U1432 ( .A(ASYNC_CMD[8]), .B(PERIOD_CMD[8]), .S(SL_PERIOD), .Y(
        SL_CRC16[8]) );
    zbfb U1433 ( .A(SL_CRC16[9]), .Y(SL_MAXLEN[1]) );
    zmux21hb U1434 ( .A(ASYNC_CMD[9]), .B(PERIOD_CMD[9]), .S(n3613), .Y(
        SL_CRC16[9]) );
    zbfb U1435 ( .A(SL_CRC16[10]), .Y(SL_MAXLEN[2]) );
    zmux21hb U1436 ( .A(ASYNC_CMD[10]), .B(PERIOD_CMD[10]), .S(n3613), .Y(
        SL_CRC16[10]) );
    zbfb U1437 ( .A(SL_CRC16[11]), .Y(SL_MAXLEN[3]) );
    zmux21hb U1438 ( .A(ASYNC_CMD[11]), .B(PERIOD_CMD[11]), .S(n3613), .Y(
        SL_CRC16[11]) );
    zbfb U1439 ( .A(SL_CRC16[12]), .Y(SL_MAXLEN[4]) );
    zmux21hb U1440 ( .A(ASYNC_CMD[12]), .B(PERIOD_CMD[12]), .S(SL_PERIOD), .Y(
        SL_CRC16[12]) );
    zbfb U1441 ( .A(SL_CRC16[13]), .Y(SL_MAXLEN[5]) );
    zmux21hb U1442 ( .A(ASYNC_CMD[13]), .B(PERIOD_CMD[13]), .S(n3613), .Y(
        SL_CRC16[13]) );
    zbfb U1443 ( .A(SL_CRC16[14]), .Y(SL_MAXLEN[6]) );
    zmux21hb U1444 ( .A(ASYNC_CMD[14]), .B(PERIOD_CMD[14]), .S(n3613), .Y(
        SL_CRC16[14]) );
    zbfb U1445 ( .A(SL_CRC16[15]), .Y(SL_MAXLEN[7]) );
    zmux21hb U1446 ( .A(ASYNC_CMD[15]), .B(PERIOD_CMD[15]), .S(SL_PERIOD), .Y(
        SL_CRC16[15]) );
    zor3b U1447 ( .A(PHASENXT_CMD_RXTOKEN), .B(CMDSMNXT_7), .C(CMDSMNXT_6), 
        .Y(NXTISRCV) );
    zor3b U1448 ( .A(n3384), .B(n3385), .C(n3386), .Y(CMDSMNXT_5) );
    zoai22d U1449 ( .A(PKTXEND), .B(n3387), .C(n3388), .D(n3389), .Y(
        CMDSMNXT_4) );
    zao222b U1450 ( .A(n3270), .B(n3390), .C(n3391), .D(n3392), .E(n3393), .F(
        n3269), .Y(CMDSMNXT_6) );
    zao222b U1451 ( .A(n3394), .B(n3275), .C(n3395), .D(n3390), .E(n3396), .F(
        n3391), .Y(CMDSMNXT_7) );
    zor6b U1452 ( .A(n3397), .B(n3398), .C(n3399), .D(n3400), .E(n3401), .F(
        n3402), .Y(NXTISIDL) );
    zao211b U1453 ( .A(n3271), .B(n3403), .C(n3404), .D(n3405), .Y(CMDSMNXT_12
        ) );
    zao211b U1454 ( .A(n3406), .B(n3390), .C(n3407), .D(n3408), .Y(
        PHASENXT_CMD_RXTOKEN) );
    zoai22d U1455 ( .A(PKTXEND), .B(n3409), .C(n3388), .D(n3410), .Y(
        CMDSMNXT_2) );
    zao211b U1456 ( .A(CMDSTATE_5), .B(n3418), .C(n3419), .D(n3420), .Y(
        RCV_POWERUP_COND) );
    znd8d U1457 ( .A(n3429), .B(n3430), .C(n3431), .D(n3432), .E(n3433), .F(
        n3434), .G(n3435), .H(n3436), .Y(NXTISTX) );
    zoai22d U1458 ( .A(PKTXEND), .B(n3438), .C(n3388), .D(n3439), .Y(
        CMDSMNXT_3) );
    zan4b U1459 ( .A(RXOUT), .B(SL_SP_ET_0), .C(n3442), .D(SL_TXDATASEL[0]), 
        .Y(n3441) );
    zoa21d U1460 ( .A(n3443), .B(n3444), .C(ASKREPLY), .Y(SEQERR) );
    zor6b U1461 ( .A(CMDSTATE_10), .B(n3445), .C(RCV_POWERUP_COND), .D(
        MAC_SLAVE_ACT), .E(DISPDRCV), .F(NXTISRCV), .Y(RCV_POWERUP2134) );
    zan2d U1462 ( .A(n3278), .B(n3449), .Y(SL_FORCE_CRC) );
    zan2d U1463 ( .A(n3278), .B(n3450), .Y(SL_FORCE_STUFF) );
    zor3b U1464 ( .A(TX_PERIOD_P), .B(TURNCNT_EN), .C(PKTXEND), .Y(TX_PERIOD)
         );
    zan2d U1465 ( .A(n3278), .B(n3456), .Y(SL_FORCE_PID) );
    zoa21d U1466 ( .A(n2356), .B(TXTMOUT), .C(CMDSTATE_13), .Y(TXTMOUT2366) );
    zoa21d U1467 ( .A(TXDELAY), .B(n2478), .C(CMDSTATE_14), .Y(TXDELAY2488) );
    zan3d U1468 ( .A(n3461), .B(n3462), .C(n3463), .Y(n3460) );
    zan4b U1469 ( .A(n3467), .B(n3468), .C(CMDSTATE_11), .D(n3469), .Y(n3407)
         );
    zan4b U1470 ( .A(MAC_CMDSTART), .B(n3411), .C(MAC_SLAVE_ACT), .D(n3470), 
        .Y(n3408) );
    zoa21d U1471 ( .A(RXDATA), .B(n3476), .C(n3424), .Y(n3475) );
    zan4b U1472 ( .A(n3410), .B(n3389), .C(n3439), .D(n3484), .Y(n3483) );
    zoa21d U1473 ( .A(n3426), .B(n3421), .C(EOF2), .Y(n3489) );
    zoa21d U1474 ( .A(RXDATA), .B(n3476), .C(n3492), .Y(n3491) );
    zan4b U1475 ( .A(n3269), .B(n3493), .C(n3494), .D(n3495), .Y(n3386) );
    zcx8d U1476 ( .A(n3403), .B(n3500), .C(MAC_CMDSTART), .D(n3440), .E(n3499), 
        .Y(n3498) );
    zan4b U1477 ( .A(RXDATA), .B(n3501), .C(NORMPKT), .D(n3424), .Y(n3404) );
    zoa21d U1478 ( .A(n3276), .B(n3263), .C(n3394), .Y(n3405) );
    zan4b U1479 ( .A(n3502), .B(n3503), .C(n3504), .D(n3505), .Y(n3446) );
    zoa21d U1480 ( .A(DAT0), .B(TEST_PACKET_T), .C(CMDSTATE_5), .Y(n3457) );
    zoa21d U1481 ( .A(n3510), .B(n3511), .C(n3277), .Y(n3458) );
    zoa21d U1482 ( .A(n3512), .B(n3513), .C(n3277), .Y(n3448) );
    zoa21d U1483 ( .A(RXTOKENPHASE), .B(CMDSTATE_6), .C(RXDATA), .Y(n3443) );
    zoa21d U1484 ( .A(RXTOKENPHASE), .B(DATAIN), .C(RXACK), .Y(n3444) );
    zoa21d U1485 ( .A(n3275), .B(n3481), .C(CMDSTATE_10), .Y(n3515) );
    zmux21ld U1486 ( .A(ASYNC_CMD[29]), .B(PERIOD_CMD[29]), .S(n3613), .Y(
        n3463) );
    zmux21ld U1487 ( .A(ASYNC_CMD[30]), .B(PERIOD_CMD[30]), .S(n3613), .Y(
        n3462) );
    zmux21ld U1488 ( .A(ASYNC_CMD[28]), .B(PERIOD_CMD[28]), .S(n3613), .Y(
        n3461) );
    zmux21ld U1489 ( .A(ASYNC_CMD[26]), .B(PERIOD_CMD[26]), .S(n3613), .Y(
        n3519) );
    zmux21ld U1490 ( .A(ASYNC_CMD[25]), .B(PERIOD_CMD[25]), .S(n3613), .Y(
        n3520) );
    zmux21ld U1491 ( .A(ASYNC_CMD[24]), .B(PERIOD_CMD[24]), .S(n3613), .Y(
        n3521) );
    zor4b U1492 ( .A(CMDSTATE_14), .B(CMDSTATE_15), .C(n3522), .D(n3523), .Y(
        n3526) );
    zor3b U1493 ( .A(CMDSTATE_10), .B(n3526), .C(n3452), .Y(n3527) );
    zor3b U1494 ( .A(CMDSTATE_15), .B(n3522), .C(n3531), .Y(n3532) );
    zor3b U1495 ( .A(CMDSTATE_5), .B(n3523), .C(n3532), .Y(n3533) );
    zor4b U1496 ( .A(TXSOF), .B(n3517), .C(n3534), .D(n3533), .Y(n3409) );
    zor3b U1497 ( .A(CMDSTATE_0), .B(n3452), .C(n3532), .Y(n3540) );
    zor2d U1498 ( .A(n3544), .B(n3539), .Y(n3494) );
    zor3b U1499 ( .A(n3545), .B(n3526), .C(CURISTX), .Y(n3546) );
    zor3b U1500 ( .A(CMDSTATE_6), .B(n3549), .C(n3540), .Y(n3550) );
    zor4b U1501 ( .A(CMDSTATE_15), .B(n3523), .C(CMDSTATE_10), .D(CURISTX), 
        .Y(n3551) );
    zor4b U1502 ( .A(n3502), .B(n3445), .C(n3452), .D(n3532), .Y(n3553) );
    zor4b U1503 ( .A(MAC_SLAVE_ACT), .B(TEST_PACKET), .C(n3553), .D(n3412), 
        .Y(n3554) );
    zor3b U1504 ( .A(n3555), .B(n3529), .C(n3527), .Y(n3500) );
    zor3b U1505 ( .A(n3522), .B(n3468), .C(n3551), .Y(n3561) );
    zor4b U1506 ( .A(CMDSTATE_14), .B(CMDSTATE_11), .C(n3467), .D(n3551), .Y(
        n3562) );
    zor2d U1507 ( .A(n3563), .B(n3542), .Y(n3418) );
    zor4b U1508 ( .A(TXIN), .B(n3517), .C(n3564), .D(n3533), .Y(n3565) );
    zor3b U1509 ( .A(EOF1), .B(n3550), .C(n3390), .Y(n3568) );
    zor4b U1510 ( .A(TXOUT), .B(n3524), .C(n3536), .D(n3533), .Y(n3387) );
    zor4b U1511 ( .A(TXSETUP), .B(n3524), .C(n3537), .D(n3533), .Y(n3438) );
    zor3b U1512 ( .A(n3390), .B(n3573), .C(n3572), .Y(n3574) );
    zor6b U1513 ( .A(n3520), .B(SL_PID[2]), .C(n3521), .D(n3578), .E(
        SL_RXSPLIT), .F(n3273), .Y(n3577) );
    zoai22d U1514 ( .A(PERIOD_CMD[31]), .B(n3615), .C(n3460), .D(n3542), .Y(
        n3578) );
    zor4b U1515 ( .A(n3480), .B(n3483), .C(n3486), .D(n3489), .Y(n3604) );
    zao211b U1516 ( .A(n3569), .B(n3570), .C(n3605), .D(n3604), .Y(n3402) );
    zao222b U1517 ( .A(TXOUT), .B(TXSETUP), .C(TXSOF), .D(TXIN), .E(DATAIN), 
        .F(CMDSTATE_6), .Y(n3398) );
    zoa22d U1518 ( .A(n3610), .B(n3572), .C(n3390), .D(n3549), .Y(n3505) );
    zor3b U1519 ( .A(TXPING), .B(TXIN), .C(n3515), .Y(n3420) );
    zao211b U1520 ( .A(n3516), .B(n3497), .C(n3268), .D(n3464), .Y(n3392) );
    zor5b U1521 ( .A(SL_PID[1]), .B(SL_PID[0]), .C(SL_PID[3]), .D(n3519), .E(
        n3542), .Y(n3593) );
    zor5b U1522 ( .A(n3437), .B(n3268), .C(n3465), .D(n3269), .E(n3497), .Y(
        n3417) );
    zor3b U1523 ( .A(n3568), .B(n3491), .C(n3559), .Y(n3612) );
    zivh U1524 ( .A(NXTISTX), .Y(n3610) );
    zor4b U1525 ( .A(n3584), .B(n3585), .C(n3582), .D(n3583), .Y(n3514) );
    zor3b U1526 ( .A(NORMPKT), .B(TXTMOUT_EN), .C(n3558), .Y(n3592) );
    zmux21ld U1527 ( .A(ASYNC_CMD[21]), .B(PERIOD_CMD[21]), .S(SL_PERIOD), .Y(
        n3595) );
    zivh U1528 ( .A(n3595), .Y(SL_TXDATASEL[1]) );
    zor3b U1529 ( .A(n3541), .B(n3390), .C(n3577), .Y(n3598) );
endmodule


module HS_BUSTIMER ( TMOUT_PARM, W4REPLY, TMOUT, RXACTIVE, CLK60M, STSRST_, 
    ATPG_ENI );
input  [7:0] TMOUT_PARM;
input  W4REPLY, RXACTIVE, CLK60M, STSRST_, ATPG_ENI;
output TMOUT;
    wire TMCNT113_0, SPAREO6, TMCNT_2, TMCNT105_2, SPAREO0_, SPAREO8, 
        TMCNT105_5, TMCNT_EN, TMCNT_5, SPAREO1, TMCNT113_7, TMCNT_4, SPAREO9, 
        TMCNT105_4, TMCNT113_6, SPAREO0, SPAREO7, TMCNT113_1, TMCNT105_3, 
        TMCNT_3, TMCNT113_3, SPAREO5, TMCNT_1, TMCNT105_1, TMCNT105_6, TMCNT_6, 
        TMCNT_EN57, TMOUT170, SPAREO2, n156, TMCNT113_4, TMCNT_7, TMCNT105_7, 
        TMCNT113_5, SPAREO3, SPAREO1_, SPAREO4, TMCNT113_2, TMCNT105_0, 
        TMCNT_0, n220, add_39_carry_6, add_39_carry_7, add_39_carry_2, 
        add_39_carry_5, add_39_carry_4, add_39_carry_3, n221, n222, n223, n224, 
        n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
        n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
        n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
        n261, n262, n263, n264, n265;
    zoai21b SPARE615 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE612 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zaoi211b SPARE613 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zoai21b SPARE614 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    znr3b SPARE616 ( .A(SPAREO2), .B(TMCNT_EN), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE618 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE611 ( .CK(CLK60M), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zdffrb SPARE610 ( .CK(CLK60M), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE619 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb SPARE617 ( .A(SPAREO4), .Y(SPAREO5) );
    znd2b U67 ( .A(TMCNT_1), .B(n255), .Y(n228) );
    znr2b U68 ( .A(TMCNT_0), .B(n240), .Y(n235) );
    zivb U69 ( .A(TMOUT_PARM[0]), .Y(n240) );
    znr2b U70 ( .A(TMCNT_2), .B(n257), .Y(n258) );
    zivb U71 ( .A(TMOUT_PARM[2]), .Y(n257) );
    znr2b U72 ( .A(TMCNT_1), .B(n255), .Y(n256) );
    zivb U73 ( .A(TMOUT_PARM[1]), .Y(n255) );
    znd2b U74 ( .A(n234), .B(n227), .Y(n226) );
    znr2b U75 ( .A(n256), .B(n258), .Y(n234) );
    znd2b U76 ( .A(n235), .B(n228), .Y(n227) );
    znr2b U77 ( .A(n260), .B(n254), .Y(n233) );
    znr2b U78 ( .A(TMOUT_PARM[2]), .B(n259), .Y(n260) );
    znr2b U79 ( .A(TMOUT_PARM[3]), .B(n253), .Y(n254) );
    znr2b U80 ( .A(TMCNT_4), .B(n249), .Y(n250) );
    zivb U81 ( .A(TMOUT_PARM[4]), .Y(n249) );
    znr2b U82 ( .A(TMCNT_3), .B(n247), .Y(n248) );
    zivb U83 ( .A(TMOUT_PARM[3]), .Y(n247) );
    znd2b U84 ( .A(n232), .B(n225), .Y(n224) );
    znr2b U85 ( .A(n248), .B(n250), .Y(n232) );
    znd2b U86 ( .A(n233), .B(n226), .Y(n225) );
    znr2b U87 ( .A(n252), .B(n246), .Y(n231) );
    znr2b U88 ( .A(TMOUT_PARM[4]), .B(n251), .Y(n252) );
    znr2b U89 ( .A(TMOUT_PARM[5]), .B(n245), .Y(n246) );
    znr2b U90 ( .A(TMCNT_5), .B(n243), .Y(n244) );
    zivb U91 ( .A(TMOUT_PARM[5]), .Y(n243) );
    znr2b U92 ( .A(TMCNT_6), .B(n241), .Y(n242) );
    znd2b U93 ( .A(TMCNT_6), .B(n241), .Y(n237) );
    zivb U94 ( .A(TMOUT_PARM[6]), .Y(n241) );
    znd2b U95 ( .A(n230), .B(n223), .Y(n238) );
    znr2b U96 ( .A(n242), .B(n244), .Y(n230) );
    znd2b U97 ( .A(n231), .B(n224), .Y(n223) );
    znd2b U98 ( .A(n221), .B(n229), .Y(n261) );
    znd2b U99 ( .A(n222), .B(n236), .Y(n221) );
    zivb U100 ( .A(TMOUT_PARM[7]), .Y(n229) );
    znd2b U101 ( .A(TMCNT_7), .B(n239), .Y(n262) );
    znd2b U102 ( .A(n238), .B(n237), .Y(n239) );
    zivb U103 ( .A(n239), .Y(n222) );
    zan2b U104 ( .A(TMCNT105_7), .B(TMCNT_EN), .Y(TMCNT113_7) );
    zxo2b U105 ( .A(add_39_carry_7), .B(TMCNT_7), .Y(TMCNT105_7) );
    zan2b U106 ( .A(TMCNT105_6), .B(TMCNT_EN), .Y(TMCNT113_6) );
    zhadrb add_39_U1_1_6 ( .A(TMCNT_6), .B(add_39_carry_6), .CO(add_39_carry_7
        ), .S(TMCNT105_6) );
    zan2b U107 ( .A(TMCNT105_5), .B(TMCNT_EN), .Y(TMCNT113_5) );
    zhadrb add_39_U1_1_5 ( .A(TMCNT_5), .B(add_39_carry_5), .CO(add_39_carry_6
        ), .S(TMCNT105_5) );
    zan2b U108 ( .A(TMCNT105_4), .B(TMCNT_EN), .Y(TMCNT113_4) );
    zhadrb add_39_U1_1_4 ( .A(TMCNT_4), .B(add_39_carry_4), .CO(add_39_carry_5
        ), .S(TMCNT105_4) );
    zan2b U109 ( .A(TMCNT105_3), .B(TMCNT_EN), .Y(TMCNT113_3) );
    zhadrb add_39_U1_1_3 ( .A(TMCNT_3), .B(add_39_carry_3), .CO(add_39_carry_4
        ), .S(TMCNT105_3) );
    zan2b U110 ( .A(TMCNT105_2), .B(TMCNT_EN), .Y(TMCNT113_2) );
    zhadrb add_39_U1_1_2 ( .A(TMCNT_2), .B(add_39_carry_2), .CO(add_39_carry_3
        ), .S(TMCNT105_2) );
    zan2b U111 ( .A(TMCNT105_1), .B(TMCNT_EN), .Y(TMCNT113_1) );
    zhadrb add_39_U1_1_1 ( .A(TMCNT_1), .B(TMCNT_0), .CO(add_39_carry_2), .S(
        TMCNT105_1) );
    zan2b U112 ( .A(TMCNT105_0), .B(TMCNT_EN), .Y(TMCNT113_0) );
    zor2b U113 ( .A(n264), .B(W4REPLY), .Y(TMCNT_EN57) );
    znr2b U114 ( .A(RXACTIVE), .B(n265), .Y(n264) );
    zor2b U115 ( .A(n156), .B(TMOUT), .Y(TMOUT170) );
    znd2b U116 ( .A(n262), .B(n261), .Y(n156) );
    zdffqrb TMCNT_reg_7 ( .CK(CLK60M), .D(TMCNT113_7), .R(STSRST_), .Q(TMCNT_7
        ) );
    zivb U117 ( .A(TMCNT_7), .Y(n236) );
    zdffqrb TMCNT_reg_6 ( .CK(CLK60M), .D(TMCNT113_6), .R(STSRST_), .Q(TMCNT_6
        ) );
    zdffqrb TMCNT_reg_5 ( .CK(CLK60M), .D(TMCNT113_5), .R(STSRST_), .Q(TMCNT_5
        ) );
    zivb U118 ( .A(TMCNT_5), .Y(n245) );
    zdffqrb TMCNT_reg_4 ( .CK(CLK60M), .D(TMCNT113_4), .R(STSRST_), .Q(TMCNT_4
        ) );
    zivb U119 ( .A(TMCNT_4), .Y(n251) );
    zdffqrb TMCNT_reg_3 ( .CK(CLK60M), .D(TMCNT113_3), .R(STSRST_), .Q(TMCNT_3
        ) );
    zivb U120 ( .A(TMCNT_3), .Y(n253) );
    zdffqrb TMCNT_reg_2 ( .CK(CLK60M), .D(TMCNT113_2), .R(STSRST_), .Q(TMCNT_2
        ) );
    zivb U121 ( .A(TMCNT_2), .Y(n259) );
    zdffqrb TMCNT_reg_1 ( .CK(CLK60M), .D(TMCNT113_1), .R(STSRST_), .Q(TMCNT_1
        ) );
    zdffqrb TMCNT_reg_0 ( .CK(CLK60M), .D(TMCNT113_0), .R(STSRST_), .Q(TMCNT_0
        ) );
    zivb U122 ( .A(TMCNT_0), .Y(TMCNT105_0) );
    zdffqrb TMCNT_EN_reg ( .CK(CLK60M), .D(TMCNT_EN57), .R(n220), .Q(TMCNT_EN)
         );
    zivb U123 ( .A(TMCNT_EN), .Y(n265) );
    zdffqrb TMOUT_reg ( .CK(CLK60M), .D(TMOUT170), .R(STSRST_), .Q(TMOUT) );
    zivb U124 ( .A(TMOUT), .Y(n263) );
    zao21b U125 ( .A(STSRST_), .B(n263), .C(ATPG_ENI), .Y(n220) );
endmodule


module DBG_PID_MUX ( DBG_TOKEN, DBG_SENDPID, HS_TXPID, TX_PID, DBG_SEL, 
    EN_DBG_PORT, TXIN, TXOUT, TXDATA0, TXSOF, DBG_PORT_BLOCKING, CLK60M );
input  [7:0] DBG_TOKEN;
input  [7:0] DBG_SENDPID;
output [7:0] TX_PID;
input  [7:0] HS_TXPID;
input  DBG_SEL, EN_DBG_PORT, TXIN, TXOUT, TXDATA0, TXSOF, CLK60M;
output DBG_PORT_BLOCKING;
    wire TXSOF_2T, TXSOF_T, n173, n174, n175, n176, n177, n178, n179, n180;
    zor2b U32 ( .A(TXIN), .B(TXOUT), .Y(n179) );
    znd2b U33 ( .A(DBG_SEL), .B(EN_DBG_PORT), .Y(n177) );
    znr4b U34 ( .A(TXSOF_2T), .B(TXSOF), .C(TXSOF_T), .D(n175), .Y(
        DBG_PORT_BLOCKING) );
    zivb U35 ( .A(DBG_SEL), .Y(n175) );
    zao21b U36 ( .A(n178), .B(n180), .C(n177), .Y(n176) );
    zivb U37 ( .A(n179), .Y(n178) );
    zivb U38 ( .A(TXDATA0), .Y(n180) );
    zdffqb TXSOF_2T_reg ( .CK(CLK60M), .D(TXSOF_T), .Q(TXSOF_2T) );
    zdffqb TXSOF_T_reg ( .CK(CLK60M), .D(TXSOF), .Q(TXSOF_T) );
    znr3b U39 ( .A(n180), .B(n179), .C(n177), .Y(n173) );
    znr2b U40 ( .A(n178), .B(n177), .Y(n174) );
    zao222b U41 ( .A(HS_TXPID[7]), .B(n176), .C(DBG_TOKEN[7]), .D(n174), .E(
        DBG_SENDPID[7]), .F(n173), .Y(TX_PID[7]) );
    zao222b U42 ( .A(HS_TXPID[6]), .B(n176), .C(DBG_TOKEN[6]), .D(n174), .E(
        DBG_SENDPID[6]), .F(n173), .Y(TX_PID[6]) );
    zao222b U43 ( .A(HS_TXPID[5]), .B(n176), .C(DBG_TOKEN[5]), .D(n174), .E(
        DBG_SENDPID[5]), .F(n173), .Y(TX_PID[5]) );
    zao222b U44 ( .A(HS_TXPID[4]), .B(n176), .C(DBG_TOKEN[4]), .D(n174), .E(
        DBG_SENDPID[4]), .F(n173), .Y(TX_PID[4]) );
    zao222b U45 ( .A(HS_TXPID[3]), .B(n176), .C(DBG_TOKEN[3]), .D(n174), .E(
        DBG_SENDPID[3]), .F(n173), .Y(TX_PID[3]) );
    zao222b U46 ( .A(HS_TXPID[2]), .B(n176), .C(DBG_TOKEN[2]), .D(n174), .E(
        DBG_SENDPID[2]), .F(n173), .Y(TX_PID[2]) );
    zao222b U47 ( .A(HS_TXPID[1]), .B(n176), .C(DBG_TOKEN[1]), .D(n174), .E(
        DBG_SENDPID[1]), .F(n173), .Y(TX_PID[1]) );
    zao222b U48 ( .A(HS_TXPID[0]), .B(n176), .C(DBG_TOKEN[0]), .D(n174), .E(
        DBG_SENDPID[0]), .F(n173), .Y(TX_PID[0]) );
endmodule

// HS MAC

module HS_MAC ( DATA_TX, TXVALID, TXREADY, CLK60M, HRST_, HCRESET, TRST_,
		DIS_STUFF, MAXLEN, HOSTDAT, USBPOP,
		DATA_RX, RXACTIVE, RXVALID, USBDAT, RXEOPERR, RXSTUFFERR,
		/*PHYRXERR,*/ DISCHKEOPERR, PHYERR, LATCHDAT, //SLAVEMODE,
		TXADDR, TXENDP, SOFV, HUBADDR, HUBPORT, SP_SC, SP_S, SP_E,
		SP_ET, EOF1, EOF2, TD_IN, TD_OUT, TD_SETUP, TD_SPLIT, TD_PING,
		CMDSTART, SOFGEN, ISO, ASKREPLY, BABBLE, MAC_EOT, TXSOF,
		EOFTERM, DAT0, DAT1, DAT2, DATM, TMOUT_PARM, CRCERR,
		ACTLEN, PIDERR, RXNAK, RXNYET, RXSTALL, RXACK, RXDATA0,
		RXDATA1, RXDATA2, RXMDATA, RXPIDERR, TMOUT, TOGMATCH,
		RXPID, SPD, RXBCNT,
		LIGHTRST, ENISOHANDCHK, EHCIEXE, //TEST_J, TEST_K, TEST_PACKET,
		SLAVE_ACT, PERIOD_CMD, ASYNC_CMD, SL_PERIOD,
		SL_DATA_PIDERR, SL_ET_ERR, SL_SE_ERR, SL_ACK_ERR, EXEITD,
		SOF_DISCONN_CHK, SOF_DISCONN, TEST_EYE_EN,
		PTstCtrl_A_3, PTstCtrl_A_2, PTstCtrl_A_1, PTstCtrl_A_0,
        	PTstCtrl_B_3, PTstCtrl_B_2, PTstCtrl_B_1, PTstCtrl_B_0,
        	PTstCtrl_C_3, PTstCtrl_C_2, PTstCtrl_C_1, PTstCtrl_C_0,
        	PTstCtrl_D_3, PTstCtrl_D_2, PTstCtrl_D_1, PTstCtrl_D_0,
        	PTstCtrl_E_3, PTstCtrl_E_2, PTstCtrl_E_1, PTstCtrl_E_0,
        	PTstCtrl_F_3, PTstCtrl_F_2, PTstCtrl_F_1, PTstCtrl_F_0,
		PTstCtrl_G_3, PTstCtrl_G_2, PTstCtrl_G_1, PTstCtrl_G_0,
		PTstCtrl_H_3, PTstCtrl_H_2, PTstCtrl_H_1, PTstCtrl_H_0,
		TEST_J, TEST_K, TEST_PACKET, TEST_FORCE_ENABLE, TEST_EYE,
		UTM_SOF, BABOPT, FBABBLE, DISPDRCV, RCV_POWERUP,
		TXTMOUT_EN, TXDELAY_EN, TXDELAY_PARM, TURN_PARM, UTM_RUN,
		FORCE_CRCERR, DIS_NARROW_SOF, EN_CHKTOGCRC, EN_UTM_RESET,
		DBG_TOKEN, DBG_SENDPID, DBG_SEL, EN_DBG_PORT, DBG_PORT_BLOCKING,
		EN_REF_RVLD, RVLD, EN_UTM_SPDUP, TX_PERIOD,
		HS_MAC_TX_CLK60M, HS_MAC_RX_CLK60M,
		ATPG_ENI, HS_TRST_
	      );
input	HS_MAC_TX_CLK60M, HS_MAC_RX_CLK60M;
output	TX_PERIOD;
input	EN_REF_RVLD, RVLD, EN_UTM_SPDUP;
input	[7:0]	DBG_TOKEN, DBG_SENDPID;
input	DBG_SEL, EN_DBG_PORT;
output	DBG_PORT_BLOCKING;
input	EN_UTM_RESET;		// enable UTM reset if UTM hang
input	EN_CHKTOGCRC;		// enable check CRCERR even TOG mismatch
input	UTM_RUN, FORCE_CRCERR, DIS_NARROW_SOF;
input	LIGHTRST, ATPG_ENI;
output	[7:0]	DATA_TX;
output  TXVALID, TRST_;
input   TXREADY, CLK60M, HRST_, HCRESET;
input   [10:0]  SOFV;
input   [10:0]  MAXLEN;
input   [7:0]   HOSTDAT;
output  USBPOP, DIS_STUFF;
input   [7:0]   DATA_RX;
input   RXACTIVE, RXVALID;
output  [7:0]   USBDAT;
input   [6:0]   TXADDR;
input   [3:0]   TXENDP;
input   [6:0]   HUBADDR, HUBPORT;
input   [1:0]   SP_ET;
input   SP_SC, SP_S, SP_E;
input   RXEOPERR, RXSTUFFERR, /*PHYRXERR,*/ DISCHKEOPERR;
output  LATCHDAT, PHYERR, ASKREPLY, BABBLE;
input	EOF1, EOF2, TD_IN, TD_OUT, TD_SETUP, TD_SPLIT, //SLAVEMODE,
	CMDSTART, SOFGEN, ISO, DAT0, DAT1, DAT2, DATM;
input	[7:0]	TMOUT_PARM;	// parameter for timeout
output	MAC_EOT, TXSOF, EOFTERM, CRCERR, PIDERR;
output	[10:0]	ACTLEN, RXBCNT;
output	RXNAK, RXNYET, RXSTALL, RXACK, TMOUT;
output	RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXPIDERR;
output	[7:0]	RXPID;
input	TD_PING;
output	TOGMATCH, SPD;
input	ENISOHANDCHK;	// check RXHAND in ISO transaction or not
input	EHCIEXE;	// EHCI control start processing TDs
output	TEST_J, TEST_K;	// test J/K state
output	TEST_PACKET;	// test_packet state
output	TEST_EYE;	// test eye pattern
input	SLAVE_ACT;	// slave mode is activated
input	[31:0]	PERIOD_CMD;	// periodic response command in slave mode
input	[31:0]	ASYNC_CMD;	// async response command in slave mode
output	SL_PERIOD;	// execute periodic command in slave mode
output	SL_DATA_PIDERR, SL_ET_ERR, SL_SE_ERR, SL_ACK_ERR;
input	EXEITD;		// iTD needs to check DATA PID sequence
input	SOF_DISCONN_CHK, TEST_EYE_EN;
output	SOF_DISCONN;
input	PTstCtrl_A_3, PTstCtrl_A_2, PTstCtrl_A_1, PTstCtrl_A_0,
       	PTstCtrl_B_3, PTstCtrl_B_2, PTstCtrl_B_1, PTstCtrl_B_0,
       	PTstCtrl_C_3, PTstCtrl_C_2, PTstCtrl_C_1, PTstCtrl_C_0,
       	PTstCtrl_D_3, PTstCtrl_D_2, PTstCtrl_D_1, PTstCtrl_D_0,
        PTstCtrl_E_3, PTstCtrl_E_2, PTstCtrl_E_1, PTstCtrl_E_0,
        PTstCtrl_F_3, PTstCtrl_F_2, PTstCtrl_F_1, PTstCtrl_F_0,
	PTstCtrl_G_3, PTstCtrl_G_2, PTstCtrl_G_1, PTstCtrl_G_0,
        PTstCtrl_H_3, PTstCtrl_H_2, PTstCtrl_H_1, PTstCtrl_H_0;
output	/*TEST_J, TEST_K, TEST_PACKET,*/ TEST_FORCE_ENABLE, UTM_SOF;
input	BABOPT;
output	FBABBLE;
input   DISPDRCV, TXTMOUT_EN;
output  RCV_POWERUP;
input	TXDELAY_EN;
input	[7:0]	TXDELAY_PARM;
input	[3:0]	TURN_PARM;
input	HS_TRST_;

wire [7:0] TX_PID, HS_TXPID;
wire [7:0] RXPID;
wire [15:0] CRC;
wire [7:0] RXCRCDAT, TXCRCDAT, CRCDATIN;
wire [18:0] ADRENDPS;
wire [7:0] TMOUT_PARM;
wire [10:0] RXBCNT, TXBCNT;
wire [23:0] RXADDRF;
wire [3:0] SL_PID;
wire [15:0] SL_CRC16;
wire [2:0] SL_TXDATASEL;
wire [7:0] SL_TXFIXDATA;
wire [10:0] MAXLEN, SL_MAXLEN, MAC_MAXLEN;
wire GND=1'b0;

zao21d DNT_CRCERR ( .A(EN_UTM_RESET), .B(PHYERR), .C(MAC_CRCERR), .Y(CRCERR) );

HS_MACCTL HS_MACCTL ( .NEWCMD(NEWCMD), .EOF1(T_EOF1), .EOF2(T_EOF2),
	.TD_IN(TD_IN), .TD_OUT(TD_OUT), .TD_SETUP(TD_SETUP),
	.TD_SPLIT(TD_SPLIT), .MAC_CMDSTART(MAC_CMDSTART), .SOFGEN(SOFGEN),
	//.CLK60M(CLK60M), .ASKREPLY(ASKREPLY), .ISO(ISO), .TXSPLIT(TXSPLIT),
	.CLK60M(CLK60M), .ASKREPLY(MAC_ASKREPLY), .ISO(ISO), .TXSPLIT(TXSPLIT),
	.TXACK(TXACK), .TXDATA0(TXDATA0), .TXDATA1(TXDATA1),
	.TXDATA2(TXDATA2), .TXMDATA(TXMDATA), .TXIN(TXIN), .TXOUT(TXOUT),
	.TXSOF(TXSOF), .TXSETUP(TXSETUP), .TRST_(HS_TRST_), .TXSTART(TXSTART),
	.PKTXEND(PKTXEND), .PKRVEND(PKRVEND), .RXDATA(RXDATA),
	.NORMPKT(NORMPKT), .SEQERR(SEQERR), .W4REPLY(W4REPLY), .RXACK(RXACK),
	.MAC_EOT(MAC_EOT), .EOFTERM(EOFTERM),
	.DAT0(DAT0), .DAT1(DAT1), .DAT2(DAT2), .DATM(DATM),
	//.RXDATA0(RXDATA0), .RXDATA1(RXDATA1), .RXDATA2(RXDATA2),
	.TD_PING(TD_PING), .TXPING(TXPING), .SP_SC(SP_SC),
	.TEST_PACKET(TEST_PACKET), .MAC_SLAVE_ACT(MAC_SLAVE_ACT),
	.RXSOF(RXSOF), .RXIN(RXIN), .RXOUT(RXOUT), .RXSPLIT(RXSPLIT),
	.RXPING(RXPING), .RXSETUP(RXSETUP), .RXTOKENPHASE(RXTOKENPHASE),
	.PERIOD_CMD(PERIOD_CMD), .ASYNC_CMD(ASYNC_CMD), .RXADDRF(RXADDRF),
	.DATAIN(DATAIN), .RXPID(RXPID), .SL_TOGMATCH(SL_TOGMATCH),
	.SL_PID(SL_PID), .SL_CRC16(SL_CRC16), //.STSRST_(STSRST_),
	.SL_PERIOD(SL_PERIOD), /*.MAC_DAT0(MAC_DAT0), .MAC_DAT1(MAC_DAT1),
	.MAC_DAT2(MAC_DAT2), .MAC_DATM(MAC_DATM)*/
	.SL_TXDATASEL(SL_TXDATASEL), .SL_TXFIXDATA(SL_TXFIXDATA),
	.SL_FORCE_CRC(SL_FORCE_CRC), .SL_FORCE_PID(SL_FORCE_PID),
	.SL_FORCE_STUFF(SL_FORCE_STUFF), .SL_DATA_PIDERR(SL_DATA_PIDERR),
	.SL_ET_ERR(SL_ET_ERR), .SL_SE_ERR(SL_SE_ERR),
	.SL_ACK_ERR(SL_ACK_ERR), .SL_MAXLEN(SL_MAXLEN),
	.DISPDRCV(DISPDRCV), .RCV_POWERUP(RCV_POWERUP),
	.TXTMOUT_EN(TXTMOUT_EN), .TMOUT_PARM(TMOUT_PARM),
	.TXDELAY_EN(TXDELAY_EN), .TXDELAY_PARM(TXDELAY_PARM),
	.TURNCNT_EN(TURNCNT_EN), .TX_PERIOD(TX_PERIOD) );

HS_TXCTL HS_TXCTL ( .DATA_TX(DATA_TX), .TXVALID(TXVALID), .TXREADY(TXREADY),
	// sync TXREADY from UTM with posedge CLK60M for correcting timing
	//.TXREADY(TXREADY_SYNC),
        .CLK60M(HS_MAC_TX_CLK60M), .TXSTART(TXSTART), .STSRST_(STSRST_),
        .TX_PID(TX_PID), .CRC(CRC), .TXSOF(TXSOF),
        .TOKEN(TOKEN), .DATPKT(DATPKT), .HANDSHK(HANDSHK),
        .SPLIT(SPLIT), .TRST_(HS_TRST_), .DIS_STUFF(DIS_STUFF),
        .MAXLEN(MAC_MAXLEN), .HOSTDAT(HOSTDAT), .TXCRCEN(TXCRCEN),
        .TXCRCRST(TXCRCRST), .ADRENDPS(ADRENDPS), .USBPOP(USBPOP),
	.PKTXEND(PKTXEND), .TXCRCDAT(TXCRCDAT), .TXBCNT(TXBCNT),
	.TEST_J(TEST_J), .TEST_K(TEST_K), .SL_TXDATASEL(SL_TXDATASEL),
	.SL_TXFIXDATA(SL_TXFIXDATA), .SL_FORCE_CRC(SL_FORCE_CRC),
	.FORCE_CRCERR(FORCE_CRCERR),
	.SL_FORCE_STUFF(SL_FORCE_STUFF), .TEST_PACKET(TEST_PACKET),
	.SOF_DISCONN_CHK(SOF_DISCONN_CHK), .SOF_DISCONN(SOF_DISCONN),
	.TXCRCPHASE(TXCRCPHASE), .TEST_EYE(TEST_EYE),
	.TURN_PARM(TURN_PARM), .DIS_NARROW_SOF(DIS_NARROW_SOF),
	.EN_UTM_SPDUP(EN_UTM_SPDUP), .TURNCNT_EN(TURNCNT_EN),
	.ATPG_ENI(ATPG_ENI) );

HS_RXCTL HS_RXCTL ( .DATA_RX(DATA_RX), .RXACTIVE(RXACTIVE), .RXVALID(RXVALID),
        //.CLK60M(CLK60M), .ASKREPLY(ASKREPLY), .TRST_(HS_TRST_),
        .CLK60M(HS_MAC_RX_CLK60M), .ASKREPLY(MAC_ASKREPLY), .TRST_(HS_TRST_),
	.USBDAT(USBDAT), .PIDERR(PIDERR), .RXPID(RXPID), .RXDATA(RXDATA),
        .RXHAND(RXHAND), .RXSTUFFERR(RXSTUFFERR), .STSRST_(STSRST_),
        .LATCHDAT(LATCHDAT), .RXCRCEN(RXCRCEN), .RXCRCRST(RXCRCRST),
        .RXCRCDAT(RXCRCDAT), .LATCHPID(LATCHPID), .CRCHK(CRCHK),
	.PKRVEND(PKRVEND), .RXEOPERR(RXEOPERR), //.PHYRXERR(PHYRXERR),
	//.DISCHKEOPERR(DISCHKEOPERR), .PHYERR(PHYERR), .CRCERR(CRCERR),
	.DISCHKEOPERR(DISCHKEOPERR), .PHYERR(PHYERR), .CRCERR(MAC_CRCERR),
	.NORMPKT(NORMPKT), .EOF2(T_EOF2), .TMOUT(TMOUT), .MAXLEN(MAC_MAXLEN),
	.BABBLE(BABBLE), .RXBCNT(RXBCNT), .DAT0(DAT0),
	.DAT1(DAT1), .DAT2(DAT2), .DATM(DATM),
        .RXDATA0(RXDATA0), .RXDATA1(RXDATA1), .RXDATA2(RXDATA2),
	.RXMDATA(RXMDATA), .TOGMATCH(TOGMATCH), .SPD(SPD),
	.RXACK(RXACK), .ISO(ISO), .RXTOKENPHASE(RXTOKENPHASE),
	.RXSOF(RXSOF), .RXTOKEN(RXTOKEN), .RXADDRF(RXADDRF),
	.DATAIN(DATAIN), .MAC_SLAVE_ACT(MAC_SLAVE_ACT),
	.SL_TOGMATCH(SL_TOGMATCH), .EXEITD(EXEITD),
	.EN_CHKTOGCRC(EN_CHKTOGCRC),
	.EN_REF_RVLD(EN_REF_RVLD), .RVLD(RVLD) );

MACETC  MACETC  ( .MAC_ASKREPLY(MAC_ASKREPLY), .ASKREPLY(ASKREPLY),
		  .EN_UTM_RESET(EN_UTM_RESET),
		  .TXCRCEN(TXCRCEN), .RXCRCEN(RXCRCEN),
                  .CRCEN(CRCEN), .TXCRCDAT(TXCRCDAT), .RXCRCDAT(RXCRCDAT),
                  .CRCDATIN(CRCDATIN), .TXCRCRST(TXCRCRST),
                  .RXCRCRST(RXCRCRST), .CRCRST(CRCRST), .DATPKT(DATPKT),
                  .RXDATA(RXDATA), .CRC16(CRC16), .TXADDR(TXADDR),
                  .TXENDP(TXENDP), .TXSOF(TXSOF), .SOFV(SOFV),
                  .ADRENDPS(ADRENDPS), .HUBADDR(HUBADDR), .HUBPORT(HUBPORT),
                  .SPLIT(SPLIT), .SP_SC(SP_SC), .SP_S(SP_S), .SP_E(SP_E),
                  .SP_ET(SP_ET), .NEWCMD(NEWCMD), .TRST_(TRST_),
		  .STSRST_(STSRST_), .HRST_(HRST_), .HCRESET(HCRESET),
		  .TD_IN(TD_IN), .TXBCNT(TXBCNT), .RXBCNT(RXBCNT),
		  .ACTLEN(ACTLEN), .USBPOP(USBPOP), //.LATCHDAT(LATCHDAT),
		  .LIGHTRST(LIGHTRST), .EHCIEXE(EHCIEXE), .CLK60M(CLK60M),
		  .EOF1(EOF1), .EOF2(EOF2), .TEST_PACKET(TEST_PACKET),
		  .T_EOF1(T_EOF1), .T_EOF2(T_EOF2), .CMDSTART(CMDSTART),
		  .MAC_CMDSTART(MAC_CMDSTART), .SLAVE_ACT(SLAVE_ACT),
		  .MAC_SLAVE_ACT(MAC_SLAVE_ACT), .MAXLEN(MAXLEN),
		  .SL_MAXLEN(SL_MAXLEN), .MAC_MAXLEN(MAC_MAXLEN),
		  .PTstCtrl_A_3(PTstCtrl_A_3), .PTstCtrl_A_2(PTstCtrl_A_2),
        	  .PTstCtrl_A_1(PTstCtrl_A_1), .PTstCtrl_A_0(PTstCtrl_A_0),
        	  .PTstCtrl_B_3(PTstCtrl_B_3), .PTstCtrl_B_2(PTstCtrl_B_2),
        	  .PTstCtrl_B_1(PTstCtrl_B_1), .PTstCtrl_B_0(PTstCtrl_B_0),
        	  .PTstCtrl_C_3(PTstCtrl_C_3), .PTstCtrl_C_2(PTstCtrl_C_2),
        	  .PTstCtrl_C_1(PTstCtrl_C_1), .PTstCtrl_C_0(PTstCtrl_C_0),
        	  .PTstCtrl_D_3(PTstCtrl_D_3), .PTstCtrl_D_2(PTstCtrl_D_2),
        	  .PTstCtrl_D_1(PTstCtrl_D_1), .PTstCtrl_D_0(PTstCtrl_D_0),
        	  .PTstCtrl_E_3(PTstCtrl_E_3), .PTstCtrl_E_2(PTstCtrl_E_2),
        	  .PTstCtrl_E_1(PTstCtrl_E_1), .PTstCtrl_E_0(PTstCtrl_E_0),
        	  .PTstCtrl_F_3(PTstCtrl_F_3), .PTstCtrl_F_2(PTstCtrl_F_2),
        	  .PTstCtrl_F_1(PTstCtrl_F_1), .PTstCtrl_F_0(PTstCtrl_F_0),
		  .PTstCtrl_G_3(PTstCtrl_G_3), .PTstCtrl_G_2(PTstCtrl_G_2),
		  .PTstCtrl_G_1(PTstCtrl_G_1), .PTstCtrl_G_0(PTstCtrl_G_0),
		  .PTstCtrl_H_3(PTstCtrl_H_3), .PTstCtrl_H_2(PTstCtrl_H_2),
		  .PTstCtrl_H_1(PTstCtrl_H_1), .PTstCtrl_H_0(PTstCtrl_H_0),
		  .TEST_J(TEST_J), .TEST_K(TEST_K), .UTM_SOF(UTM_SOF),
		  .TEST_FORCE_ENABLE(TEST_FORCE_ENABLE),
		  .TXCRCPHASE(TXCRCPHASE), .TXVALID(TXVALID),
		  .RXACTIVE(RXACTIVE), .BABOPT(BABOPT), .FBABBLE(FBABBLE),
		  .TEST_EYE_EN(TEST_EYE_EN), .TEST_EYE(TEST_EYE),
		  .ATPG_ENI(ATPG_ENI), .HS_TRST_(HS_TRST_),
		  .UTM_TXREADY(TXREADY), .TXREADY_SYNC(TXREADY_SYNC),
		  .UTM_RUN(UTM_RUN) );

HS_CRC  HS_CRC ( .DATAIN(CRCDATIN), .CRC(CRC), .CRC16(CRC16),
                 .CLK60M(CLK60M), .CRCRST(CRCRST), .CRCEN(CRCEN),
                 .ADRENDPS(ADRENDPS), .SPLIT(SPLIT), .RXDATA(RXDATA),
                 //.STSRST_(STSRST_), .CRCHK(CRCHK), .CRCERR(CRCERR),
                 .STSRST_(STSRST_), .CRCHK(CRCHK), .CRCERR(MAC_CRCERR),
		 .MAC_SLAVE_ACT(MAC_SLAVE_ACT), .SL_CRC16(SL_CRC16) );

HS_PIDENC HS_PIDENC ( .TXOUT(TXOUT), .TXIN(TXIN), .TXSOF(TXSOF),
                .TXSETUP(TXSETUP), .TXDATA0(TXDATA0), .TXDATA1(TXDATA1),
                .TXDATA2(TXDATA2), .TXMDATA(TXMDATA), .TXACK(TXACK),

                //.TXNAK(TXNAK), .TXSTALL(TXSTALL), .TXNYET(TXNYET),
                //.TXERR(TXERR), .TXSPLIT(TXSPLIT), .TXPING(TXPING),
		.TXNAK(GND), .TXSTALL(GND), .TXNYET(GND),
                .TXERR(GND), .TXSPLIT(TXSPLIT), .TXPING(TXPING),

                //.TX_PID(TX_PID), .TOKEN(TOKEN), .DATPKT(DATPKT),
                .TX_PID(HS_TXPID), .TOKEN(TOKEN), .DATPKT(DATPKT),
                .HANDSHK(HANDSHK), .SPLIT(SPLIT),
		.MAC_SLAVE_ACT(MAC_SLAVE_ACT), .SL_PID(SL_PID),
		.SL_FORCE_PID(SL_FORCE_PID) );

HS_PIDEC HS_PIDEC ( .RXPID(RXPID), .RXACK(RXACK), .RXDATA0(RXDATA0),
                .RXDATA1(RXDATA1), .RXDATA2(RXDATA2), .RXMDATA(RXMDATA),
                .RXNAK(RXNAK), .RXSTALL(RXSTALL), .RXNYET(RXNYET),
                .RXERR(RXPIDERR), .RXHAND(RXHAND), .RXTOKEN(RXTOKEN),
                .PIDERR(PIDERR), .RXOUT(RXOUT), .RXIN(RXIN), .RXDATA(RXDATA),
                .RXSOF(RXSOF), .RXSETUP(RXSETUP), .RXPING(RXPING),
                .RXSPLIT(RXSPLIT), .STSRST_(STSRST_), .LATCHPID(LATCHPID),
                .ISO(ISO), .SEQERR(SEQERR), .MAC_SLAVE_ACT(MAC_SLAVE_ACT),
		.ENISOHANDCHK(ENISOHANDCHK), .ATPG_ENI(ATPG_ENI) );

HS_BUSTIMER HS_BUSTIMER ( .TMOUT_PARM(TMOUT_PARM), .W4REPLY(W4REPLY),
		.TMOUT(TMOUT), .RXACTIVE(RXACTIVE), .CLK60M(CLK60M),
		.STSRST_(STSRST_), .ATPG_ENI(ATPG_ENI) );

DBG_PID_MUX DBG_PID_MUX ( .DBG_TOKEN(DBG_TOKEN), .DBG_SENDPID(DBG_SENDPID),
		.HS_TXPID(HS_TXPID), .TX_PID(TX_PID), .DBG_SEL(DBG_SEL),
                .EN_DBG_PORT(EN_DBG_PORT), .TXIN(TXIN), .TXOUT(TXOUT),
		.TXDATA0(TXDATA0), .TXSOF(TXSOF),
		.DBG_PORT_BLOCKING(DBG_PORT_BLOCKING), .CLK60M(CLK60M) );

endmodule


module ASYNCFLOW ( ASYNC_EN, PCIEND, GEN_PERR, DWNUM, EHCIREQ, RUN, ASYNC_ACT, 
    PARSEQHEND1, PARSEQHEND2, QH_PARSE_GO1, QH_PARSE_GO2, QHPARSING1, 
    QHPARSING2, QHIDLE1, QHIDLE2, QH_ACT1, QH_ACT2, ASYNC_EXE1, ASYNC_EXE2, 
    QHCIREQ1, QHCIREQ2, QHCIGNT1, QHCIGNT2, QH_CACHE_EN1, QH_CACHE_EN2, 
    DWOFFSET, ASYNCLISTADDR, CACHE_ADDR1, CACHE_ADDR2, CACHE_SEL, 
    CACHE_INVALID1, CACHE_INVALID2, LIST_SEL, QTDEXE1, QTDEXE2, HEADSEEN1, 
    HEADSEEN2, ASYNC_EMPTY1, ASYNC_EMPTY2, RECLAMATION, EHCISLEEP, EHCIRESTART, 
    START_EVENT, NAKCNTSM, NAKCNTSMNXT, INTASYNC_EN, INTASYNC, INTDOORBELL, 
    LTINT_PCLK, INTASYNC_S, QHASYNCINT, SWDBG, RUN_C, FROZEN, QCMDSTART1, 
    QCMDSTART2, PCICLK, TRST_ );
output [3:0] DWNUM;
output [3:0] DWOFFSET;
output [26:0] CACHE_ADDR2;
output [1:0] NAKCNTSMNXT;
output [1:0] NAKCNTSM;
input  [31:0] ASYNCLISTADDR;
output [26:0] CACHE_ADDR1;
input  ASYNC_EN, PCIEND, GEN_PERR, RUN, PARSEQHEND1, PARSEQHEND2, QHPARSING1, 
    QHPARSING2, QHIDLE1, QHIDLE2, QHCIREQ1, QHCIREQ2, CACHE_INVALID1, 
    CACHE_INVALID2, LIST_SEL, QTDEXE1, QTDEXE2, HEADSEEN1, HEADSEEN2, 
    ASYNC_EMPTY1, ASYNC_EMPTY2, EHCIRESTART, INTASYNC_EN, INTASYNC, 
    INTDOORBELL, LTINT_PCLK, SWDBG, QCMDSTART1, QCMDSTART2, PCICLK, TRST_;
output EHCIREQ, ASYNC_ACT, QH_PARSE_GO1, QH_PARSE_GO2, QH_ACT1, QH_ACT2, 
    ASYNC_EXE1, ASYNC_EXE2, QHCIGNT1, QHCIGNT2, QH_CACHE_EN1, QH_CACHE_EN2, 
    CACHE_SEL, RECLAMATION, EHCISLEEP, START_EVENT, INTASYNC_S, QHASYNCINT, 
    RUN_C, FROZEN;
    wire CACHE_ADDR1721_22, CACHE_HIT, ASYNCSMNXT_4, SPAREO6, 
        CACHE_ADDR2759_15, CACHE_ADDR2759_9, CACHE_ADDR2759_20, 
        CACHE_ADDR2759_0, HEADSEEN_PRE, CACHE_ADDR1721_17, CACHE_ADDR1721_6, 
        CACHE_ADDR1721_1, CACHE_ADDR1721_10, CACHE_ADDR2759_7, SPAREO0_, 
        LIST_SEL_T, SPAREO8, QH_ACT_SEL552, CACHE_ADDR1721_19, 
        CACHE_ADDR1721_8, EHCISLEEP1231, CACHE_ADDR2759_12, ASYNCSMNXT_3, 
        SPAREO1, CACHE_ADDR1721_25, QHASYNCINT1448, EHCIRESTART_T, 
        CACHE_ADDR2759_6, CACHE_ADDR2759_26, EXE_HALT, ASYNCSM_3, 
        CACHE_ADDR1721_0, CACHE_ADDR1721_11, CACHE_ADDR1721_24, 
        CACHE_ADDR2759_13, SPAREO0, CACHE_ADDR1721_18, CACHE_ADDR1721_9, 
        QH_PARSE_GO1_T, CACHEHIT1, CACHE_ADDR2759_8, ASYNCSM_4, SPAREO7, 
        CACHE_ADDR2759_14, CACHE_ADDR1721_23, CACHE_ADDR1721_16, 
        PHASENXT_ParseQH, EXE_HALT_pre, RECLAMATION1194, CACHE_ADDR1721_7, 
        CACHE_ADDR2759_21, CACHE_ADDR2759_1, CACHE_ADDR1721_21, RUN_T, 
        CACHE_ADDR2759_16, CACHE_SEL_PRE, SPAREO5, FROZEN1366, 
        EHCIRESTART_SYNC313, DOORCNT_1, DOORCNT1410_0, HEADSEEN_2T, 
        CACHE_ADDR2759_3, CACHE_ADDR2759_23, CACHE_ADDR1721_5, 
        CACHE_ADDR1721_14, ASYNCSM_1, CACHE_ADDR1721_13, CACHE_ADDR1721_2, 
        CACHE_ADDR2759_24, CACHE_ADDR2759_4, CACHE_ADDR2759_18, HEADSEEN_T, 
        EHCIRESTART_SYNC, QH_PARSE_GO2_T, ASYNCSMNXT_0, SPAREO2, 
        CACHE_ADDR2759_11, CACHE_ADDR1721_26, CACHE_ADDR2759_19, ASYNCSM_0, 
        CACHE_ADDR2759_25, CACHE_ADDR2759_5, CACHE_ADDR1721_12, 
        CACHE_ADDR1721_3, ASYNCSMNXT_1, SPAREO3, CACHE_ADDR2759_10, SPAREO1_, 
        TRANEXED1268, CACHEHIT2, CACHE_ADDR2759_17, HEADSEEN, RUN_ASYNC, 
        PHASE_ParseQH, SPAREO4, CACHE_ADDR1721_20, CACHE_ADDR1721_4, 
        CACHE_ADDR1721_15, CACHE_ADDR2759_2, CACHE_ADDR2759_22, DOORCNT1410_1, 
        TRANEXED, DOORCNT_0, n1613, n1614, n1616, n1617, n1618, n1619, n1620, 
        n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, 
        n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, 
        n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, 
        n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, 
        n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, 
        n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, 
        n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, 
        n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, 
        n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, 
        n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, 
        n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
        n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, 
        n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, 
        n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, 
        n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, 
        n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, 
        n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, 
        n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, 
        n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, 
        n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, 
        n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830;
    assign DWNUM[3] = 1'b1;
    assign DWNUM[2] = 1'b0;
    assign DWNUM[1] = 1'b1;
    assign DWNUM[0] = 1'b1;
    assign DWOFFSET[3] = 1'b0;
    assign DWOFFSET[2] = 1'b0;
    assign DWOFFSET[1] = 1'b0;
    assign DWOFFSET[0] = 1'b0;
    znd3b SPARE839 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE830 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE837 ( .A(SPAREO4), .Y(SPAREO5) );
    znr3b SPARE836 ( .A(SPAREO2), .B(ASYNCSM_1), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE838 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE831 ( .CK(PCICLK), .D(SPAREO7), .R(TRST_), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zaoi211b SPARE833 ( .A(SPAREO4), .B(CACHEHIT2), .C(SPAREO6), .D(
        ASYNCSMNXT_1), .Y(SPAREO8) );
    zoai21b SPARE834 ( .A(SPAREO0), .B(SPAREO8), .C(START_EVENT) );
    zoai21b SPARE835 ( .A(SPAREO1), .B(EXE_HALT_pre), .C(CACHE_HIT), .Y(
        SPAREO3) );
    zaoi211b SPARE832 ( .A(SPAREO0), .B(CACHEHIT1), .C(SPAREO1_), .D(RUN_ASYNC
        ), .Y(SPAREO2) );
    zxo2b U502 ( .A(n1715), .B(ASYNCLISTADDR[25]), .Y(n1803) );
    zxo2b U503 ( .A(n1714), .B(ASYNCLISTADDR[5]), .Y(n1804) );
    zxo2b U504 ( .A(n1713), .B(ASYNCLISTADDR[13]), .Y(n1805) );
    zxo2b U505 ( .A(n1712), .B(ASYNCLISTADDR[6]), .Y(n1806) );
    zxo2b U506 ( .A(n1718), .B(ASYNCLISTADDR[11]), .Y(n1817) );
    zxo2b U507 ( .A(n1716), .B(ASYNCLISTADDR[18]), .Y(n1816) );
    zxo2b U508 ( .A(n1717), .B(ASYNCLISTADDR[24]), .Y(n1815) );
    zxo2b U509 ( .A(n1722), .B(ASYNCLISTADDR[29]), .Y(n1808) );
    zxo2b U510 ( .A(n1721), .B(ASYNCLISTADDR[17]), .Y(n1809) );
    zxo2b U511 ( .A(n1720), .B(ASYNCLISTADDR[30]), .Y(n1810) );
    zxo2b U512 ( .A(n1719), .B(ASYNCLISTADDR[10]), .Y(n1811) );
    zxo2b U513 ( .A(n1725), .B(ASYNCLISTADDR[7]), .Y(n1814) );
    zxo2b U514 ( .A(n1723), .B(ASYNCLISTADDR[26]), .Y(n1813) );
    zxo2b U515 ( .A(n1724), .B(ASYNCLISTADDR[12]), .Y(n1812) );
    zxo2b U516 ( .A(ASYNCLISTADDR[15]), .B(CACHE_ADDR1[10]), .Y(n1769) );
    zxo2b U517 ( .A(ASYNCLISTADDR[8]), .B(CACHE_ADDR1[3]), .Y(n1768) );
    zxo2b U518 ( .A(ASYNCLISTADDR[9]), .B(CACHE_ADDR1[4]), .Y(n1767) );
    zxo2b U519 ( .A(ASYNCLISTADDR[22]), .B(CACHE_ADDR1[17]), .Y(n1772) );
    zxo2b U520 ( .A(ASYNCLISTADDR[27]), .B(CACHE_ADDR1[22]), .Y(n1771) );
    zxo2b U521 ( .A(ASYNCLISTADDR[23]), .B(CACHE_ADDR1[18]), .Y(n1770) );
    zxo2b U522 ( .A(ASYNCLISTADDR[14]), .B(CACHE_ADDR1[9]), .Y(n1764) );
    zxo2b U523 ( .A(ASYNCLISTADDR[19]), .B(CACHE_ADDR1[14]), .Y(n1763) );
    zxo2b U524 ( .A(ASYNCLISTADDR[28]), .B(CACHE_ADDR1[23]), .Y(n1766) );
    zxo2b U525 ( .A(ASYNCLISTADDR[31]), .B(CACHE_ADDR1[26]), .Y(n1765) );
    zxo2b U526 ( .A(n1695), .B(ASYNCLISTADDR[24]), .Y(n1787) );
    zxo2b U527 ( .A(n1694), .B(ASYNCLISTADDR[18]), .Y(n1788) );
    zxo2b U528 ( .A(n1693), .B(ASYNCLISTADDR[19]), .Y(n1789) );
    zxo2b U529 ( .A(n1692), .B(ASYNCLISTADDR[26]), .Y(n1790) );
    zxo2b U530 ( .A(n1698), .B(ASYNCLISTADDR[8]), .Y(n1801) );
    zxo2b U531 ( .A(n1696), .B(ASYNCLISTADDR[7]), .Y(n1800) );
    zxo2b U532 ( .A(n1697), .B(ASYNCLISTADDR[23]), .Y(n1799) );
    zxo2b U533 ( .A(n1702), .B(ASYNCLISTADDR[25]), .Y(n1792) );
    zxo2b U534 ( .A(n1701), .B(ASYNCLISTADDR[31]), .Y(n1793) );
    zxo2b U535 ( .A(n1700), .B(ASYNCLISTADDR[17]), .Y(n1794) );
    zxo2b U536 ( .A(n1699), .B(ASYNCLISTADDR[22]), .Y(n1795) );
    zxo2b U537 ( .A(n1705), .B(ASYNCLISTADDR[20]), .Y(n1798) );
    zxo2b U538 ( .A(n1703), .B(ASYNCLISTADDR[9]), .Y(n1797) );
    zxo2b U539 ( .A(n1704), .B(ASYNCLISTADDR[27]), .Y(n1796) );
    zxo2b U540 ( .A(CACHE_ADDR2[5]), .B(ASYNCLISTADDR[10]), .Y(n1759) );
    zxo2b U541 ( .A(CACHE_ADDR2[0]), .B(ASYNCLISTADDR[5]), .Y(n1758) );
    zxo2b U542 ( .A(CACHE_ADDR2[1]), .B(ASYNCLISTADDR[6]), .Y(n1757) );
    zxo2b U543 ( .A(ASYNCLISTADDR[15]), .B(CACHE_ADDR2[10]), .Y(n1762) );
    zxo2b U544 ( .A(ASYNCLISTADDR[14]), .B(CACHE_ADDR2[9]), .Y(n1761) );
    zxo2b U545 ( .A(ASYNCLISTADDR[16]), .B(CACHE_ADDR2[11]), .Y(n1760) );
    zxo2b U546 ( .A(CACHE_ADDR2[24]), .B(ASYNCLISTADDR[29]), .Y(n1754) );
    zxo2b U547 ( .A(CACHE_ADDR2[25]), .B(ASYNCLISTADDR[30]), .Y(n1753) );
    zxo2b U548 ( .A(CACHE_ADDR2[16]), .B(ASYNCLISTADDR[21]), .Y(n1756) );
    zxo2b U549 ( .A(CACHE_ADDR2[23]), .B(ASYNCLISTADDR[28]), .Y(n1755) );
    zor2b U550 ( .A(QHIDLE1), .B(n1668), .Y(n1782) );
    zmux21lb U551 ( .A(n1673), .B(n1675), .S(CACHE_SEL), .Y(n1775) );
    zan2b U552 ( .A(QHIDLE2), .B(n1674), .Y(n1673) );
    zan2b U553 ( .A(QHIDLE1), .B(n1676), .Y(n1675) );
    zmux21lb U554 ( .A(n1665), .B(n1664), .S(QH_ACT2), .Y(n1778) );
    zor2b U555 ( .A(CACHE_SEL), .B(n1747), .Y(n1751) );
    zivb U556 ( .A(PARSEQHEND1), .Y(n1747) );
    zor2b U557 ( .A(n1734), .B(n1741), .Y(n1745) );
    zivb U558 ( .A(PARSEQHEND2), .Y(n1741) );
    zmux21lb U559 ( .A(n1632), .B(n1640), .S(QH_ACT2), .Y(n1667) );
    zmux21lb U560 ( .A(n1776), .B(n1777), .S(QH_ACT2), .Y(n1663) );
    zor2b U561 ( .A(QHPARSING1), .B(n1735), .Y(n1776) );
    zivb U562 ( .A(QHPARSING2), .Y(n1735) );
    zor2b U563 ( .A(QHPARSING2), .B(n1736), .Y(n1777) );
    zivb U564 ( .A(QHPARSING1), .Y(n1736) );
    zxo2b U565 ( .A(ASYNCLISTADDR[20]), .B(CACHE_ADDR1[15]), .Y(n1726) );
    zxo2b U566 ( .A(ASYNCLISTADDR[16]), .B(CACHE_ADDR1[11]), .Y(n1727) );
    zxo2b U567 ( .A(ASYNCLISTADDR[21]), .B(CACHE_ADDR1[16]), .Y(n1728) );
    znd8b U568 ( .A(n1812), .B(n1813), .C(n1814), .D(n1807), .E(n1815), .F(
        n1816), .G(n1817), .H(n1802), .Y(n1731) );
    zxo2b U569 ( .A(CACHE_ADDR2[7]), .B(ASYNCLISTADDR[12]), .Y(n1706) );
    zxo2b U570 ( .A(CACHE_ADDR2[6]), .B(ASYNCLISTADDR[11]), .Y(n1707) );
    zxo2b U571 ( .A(CACHE_ADDR2[8]), .B(ASYNCLISTADDR[13]), .Y(n1708) );
    znd8b U572 ( .A(n1796), .B(n1797), .C(n1798), .D(n1791), .E(n1799), .F(
        n1800), .G(n1801), .H(n1786), .Y(n1711) );
    zor2b U573 ( .A(ASYNC_EN), .B(n1632), .Y(n1774) );
    zmux21lb U574 ( .A(QHIDLE1), .B(n1774), .S(QHIDLE2), .Y(n1773) );
    zor2b U575 ( .A(CACHEHIT1), .B(CACHEHIT2), .Y(CACHE_HIT) );
    zivb U576 ( .A(CACHE_HIT), .Y(n1669) );
    zor2b U577 ( .A(ASYNCSM_0), .B(n1683), .Y(n1690) );
    zor2b U578 ( .A(ASYNCSM_1), .B(ASYNCSM_3), .Y(n1678) );
    zor2b U579 ( .A(HEADSEEN_T), .B(n1682), .Y(n1779) );
    zivb U580 ( .A(ASYNC_EN), .Y(n1659) );
    zao22b U581 ( .A(n1785), .B(n1739), .C(n1672), .D(n1637), .Y(n1660) );
    zxo2b U582 ( .A(n1678), .B(n1679), .Y(n1677) );
    zivb U583 ( .A(n1690), .Y(n1679) );
    zor2b U584 ( .A(ASYNCSM_4), .B(PHASE_ParseQH), .Y(n1683) );
    zan2b U585 ( .A(n1785), .B(n1739), .Y(n1784) );
    zivb U586 ( .A(n1684), .Y(n1785) );
    zxo2b U587 ( .A(n1681), .B(CACHE_SEL), .Y(n1680) );
    zivb U588 ( .A(n1783), .Y(n1826) );
    zxo2b U589 ( .A(QH_ACT1), .B(n1778), .Y(n1783) );
    zao22b U590 ( .A(n1646), .B(ASYNCLISTADDR[31]), .C(n1647), .D(CACHE_ADDR1
        [26]), .Y(CACHE_ADDR1721_26) );
    zao22b U591 ( .A(n1827), .B(ASYNCLISTADDR[30]), .C(n1828), .D(CACHE_ADDR1
        [25]), .Y(CACHE_ADDR1721_25) );
    zao22b U592 ( .A(n1646), .B(ASYNCLISTADDR[29]), .C(n1647), .D(CACHE_ADDR1
        [24]), .Y(CACHE_ADDR1721_24) );
    zao22b U593 ( .A(n1827), .B(ASYNCLISTADDR[28]), .C(n1828), .D(CACHE_ADDR1
        [23]), .Y(CACHE_ADDR1721_23) );
    zao22b U594 ( .A(n1646), .B(ASYNCLISTADDR[27]), .C(n1647), .D(CACHE_ADDR1
        [22]), .Y(CACHE_ADDR1721_22) );
    zao22b U595 ( .A(n1827), .B(ASYNCLISTADDR[26]), .C(n1828), .D(CACHE_ADDR1
        [21]), .Y(CACHE_ADDR1721_21) );
    zao22b U596 ( .A(n1827), .B(ASYNCLISTADDR[25]), .C(n1647), .D(CACHE_ADDR1
        [20]), .Y(CACHE_ADDR1721_20) );
    zao22b U597 ( .A(n1646), .B(ASYNCLISTADDR[24]), .C(n1828), .D(CACHE_ADDR1
        [19]), .Y(CACHE_ADDR1721_19) );
    zao22b U598 ( .A(n1646), .B(ASYNCLISTADDR[23]), .C(n1647), .D(CACHE_ADDR1
        [18]), .Y(CACHE_ADDR1721_18) );
    zao22b U599 ( .A(n1827), .B(ASYNCLISTADDR[22]), .C(n1828), .D(CACHE_ADDR1
        [17]), .Y(CACHE_ADDR1721_17) );
    zao22b U600 ( .A(n1827), .B(ASYNCLISTADDR[21]), .C(n1647), .D(CACHE_ADDR1
        [16]), .Y(CACHE_ADDR1721_16) );
    zao22b U601 ( .A(n1646), .B(ASYNCLISTADDR[20]), .C(n1828), .D(CACHE_ADDR1
        [15]), .Y(CACHE_ADDR1721_15) );
    zao22b U602 ( .A(n1646), .B(ASYNCLISTADDR[19]), .C(n1647), .D(CACHE_ADDR1
        [14]), .Y(CACHE_ADDR1721_14) );
    zao22b U603 ( .A(n1827), .B(ASYNCLISTADDR[18]), .C(n1828), .D(CACHE_ADDR1
        [13]), .Y(CACHE_ADDR1721_13) );
    zao22b U604 ( .A(n1646), .B(ASYNCLISTADDR[17]), .C(n1647), .D(CACHE_ADDR1
        [12]), .Y(CACHE_ADDR1721_12) );
    zao22b U605 ( .A(n1827), .B(ASYNCLISTADDR[16]), .C(n1828), .D(CACHE_ADDR1
        [11]), .Y(CACHE_ADDR1721_11) );
    zao22b U606 ( .A(n1646), .B(ASYNCLISTADDR[15]), .C(n1647), .D(CACHE_ADDR1
        [10]), .Y(CACHE_ADDR1721_10) );
    zao22b U607 ( .A(n1827), .B(ASYNCLISTADDR[14]), .C(n1828), .D(CACHE_ADDR1
        [9]), .Y(CACHE_ADDR1721_9) );
    zao22b U608 ( .A(n1646), .B(ASYNCLISTADDR[13]), .C(n1647), .D(CACHE_ADDR1
        [8]), .Y(CACHE_ADDR1721_8) );
    zao22b U609 ( .A(n1827), .B(ASYNCLISTADDR[12]), .C(n1828), .D(CACHE_ADDR1
        [7]), .Y(CACHE_ADDR1721_7) );
    zao22b U610 ( .A(n1646), .B(ASYNCLISTADDR[11]), .C(n1647), .D(CACHE_ADDR1
        [6]), .Y(CACHE_ADDR1721_6) );
    zao22b U611 ( .A(n1827), .B(ASYNCLISTADDR[10]), .C(n1828), .D(CACHE_ADDR1
        [5]), .Y(CACHE_ADDR1721_5) );
    zao22b U612 ( .A(n1827), .B(ASYNCLISTADDR[9]), .C(n1647), .D(CACHE_ADDR1
        [4]), .Y(CACHE_ADDR1721_4) );
    zao22b U613 ( .A(n1646), .B(ASYNCLISTADDR[8]), .C(n1828), .D(CACHE_ADDR1
        [3]), .Y(CACHE_ADDR1721_3) );
    zao22b U614 ( .A(n1646), .B(ASYNCLISTADDR[7]), .C(n1647), .D(CACHE_ADDR1
        [2]), .Y(CACHE_ADDR1721_2) );
    zao22b U615 ( .A(n1827), .B(ASYNCLISTADDR[6]), .C(n1828), .D(CACHE_ADDR1
        [1]), .Y(CACHE_ADDR1721_1) );
    zao22b U616 ( .A(n1646), .B(ASYNCLISTADDR[5]), .C(n1647), .D(CACHE_ADDR1
        [0]), .Y(CACHE_ADDR1721_0) );
    zivb U617 ( .A(n1752), .Y(n1646) );
    zor2b U618 ( .A(n1748), .B(n1751), .Y(n1752) );
    zivb U619 ( .A(n1749), .Y(n1647) );
    zor2b U620 ( .A(n1750), .B(n1748), .Y(n1749) );
    zivb U621 ( .A(n1751), .Y(n1750) );
    zivb U622 ( .A(n1752), .Y(n1827) );
    zivb U623 ( .A(n1749), .Y(n1828) );
    zao22b U624 ( .A(n1654), .B(ASYNCLISTADDR[31]), .C(n1655), .D(CACHE_ADDR2
        [26]), .Y(CACHE_ADDR2759_26) );
    zao22b U625 ( .A(n1829), .B(ASYNCLISTADDR[30]), .C(n1830), .D(CACHE_ADDR2
        [25]), .Y(CACHE_ADDR2759_25) );
    zao22b U626 ( .A(n1654), .B(ASYNCLISTADDR[29]), .C(n1655), .D(CACHE_ADDR2
        [24]), .Y(CACHE_ADDR2759_24) );
    zao22b U627 ( .A(n1829), .B(ASYNCLISTADDR[28]), .C(n1830), .D(CACHE_ADDR2
        [23]), .Y(CACHE_ADDR2759_23) );
    zao22b U628 ( .A(n1654), .B(ASYNCLISTADDR[27]), .C(n1655), .D(CACHE_ADDR2
        [22]), .Y(CACHE_ADDR2759_22) );
    zao22b U629 ( .A(n1829), .B(ASYNCLISTADDR[26]), .C(n1830), .D(CACHE_ADDR2
        [21]), .Y(CACHE_ADDR2759_21) );
    zao22b U630 ( .A(n1829), .B(ASYNCLISTADDR[25]), .C(n1655), .D(CACHE_ADDR2
        [20]), .Y(CACHE_ADDR2759_20) );
    zao22b U631 ( .A(n1654), .B(ASYNCLISTADDR[24]), .C(n1830), .D(CACHE_ADDR2
        [19]), .Y(CACHE_ADDR2759_19) );
    zao22b U632 ( .A(n1654), .B(ASYNCLISTADDR[23]), .C(n1655), .D(CACHE_ADDR2
        [18]), .Y(CACHE_ADDR2759_18) );
    zao22b U633 ( .A(n1829), .B(ASYNCLISTADDR[22]), .C(n1830), .D(CACHE_ADDR2
        [17]), .Y(CACHE_ADDR2759_17) );
    zao22b U634 ( .A(n1829), .B(ASYNCLISTADDR[21]), .C(n1655), .D(CACHE_ADDR2
        [16]), .Y(CACHE_ADDR2759_16) );
    zao22b U635 ( .A(n1654), .B(ASYNCLISTADDR[20]), .C(n1830), .D(CACHE_ADDR2
        [15]), .Y(CACHE_ADDR2759_15) );
    zao22b U636 ( .A(n1654), .B(ASYNCLISTADDR[19]), .C(n1655), .D(CACHE_ADDR2
        [14]), .Y(CACHE_ADDR2759_14) );
    zao22b U637 ( .A(n1829), .B(ASYNCLISTADDR[18]), .C(n1830), .D(CACHE_ADDR2
        [13]), .Y(CACHE_ADDR2759_13) );
    zao22b U638 ( .A(n1654), .B(ASYNCLISTADDR[17]), .C(n1655), .D(CACHE_ADDR2
        [12]), .Y(CACHE_ADDR2759_12) );
    zao22b U639 ( .A(n1829), .B(ASYNCLISTADDR[16]), .C(n1830), .D(CACHE_ADDR2
        [11]), .Y(CACHE_ADDR2759_11) );
    zao22b U640 ( .A(n1654), .B(ASYNCLISTADDR[15]), .C(n1655), .D(CACHE_ADDR2
        [10]), .Y(CACHE_ADDR2759_10) );
    zao22b U641 ( .A(n1829), .B(ASYNCLISTADDR[14]), .C(n1830), .D(CACHE_ADDR2
        [9]), .Y(CACHE_ADDR2759_9) );
    zao22b U642 ( .A(n1654), .B(ASYNCLISTADDR[13]), .C(n1655), .D(CACHE_ADDR2
        [8]), .Y(CACHE_ADDR2759_8) );
    zao22b U643 ( .A(n1829), .B(ASYNCLISTADDR[12]), .C(n1830), .D(CACHE_ADDR2
        [7]), .Y(CACHE_ADDR2759_7) );
    zao22b U644 ( .A(n1654), .B(ASYNCLISTADDR[11]), .C(n1655), .D(CACHE_ADDR2
        [6]), .Y(CACHE_ADDR2759_6) );
    zao22b U645 ( .A(n1829), .B(ASYNCLISTADDR[10]), .C(n1830), .D(CACHE_ADDR2
        [5]), .Y(CACHE_ADDR2759_5) );
    zao22b U646 ( .A(n1829), .B(ASYNCLISTADDR[9]), .C(n1655), .D(CACHE_ADDR2
        [4]), .Y(CACHE_ADDR2759_4) );
    zao22b U647 ( .A(n1654), .B(ASYNCLISTADDR[8]), .C(n1830), .D(CACHE_ADDR2
        [3]), .Y(CACHE_ADDR2759_3) );
    zao22b U648 ( .A(n1654), .B(ASYNCLISTADDR[7]), .C(n1655), .D(CACHE_ADDR2
        [2]), .Y(CACHE_ADDR2759_2) );
    zao22b U649 ( .A(n1829), .B(ASYNCLISTADDR[6]), .C(n1830), .D(CACHE_ADDR2
        [1]), .Y(CACHE_ADDR2759_1) );
    zao22b U650 ( .A(n1654), .B(ASYNCLISTADDR[5]), .C(n1655), .D(CACHE_ADDR2
        [0]), .Y(CACHE_ADDR2759_0) );
    zivb U651 ( .A(n1746), .Y(n1654) );
    zor2b U652 ( .A(n1742), .B(n1745), .Y(n1746) );
    zivb U653 ( .A(n1743), .Y(n1655) );
    zor2b U654 ( .A(n1744), .B(n1742), .Y(n1743) );
    zivb U655 ( .A(n1745), .Y(n1744) );
    zivb U656 ( .A(n1746), .Y(n1829) );
    zivb U657 ( .A(n1743), .Y(n1830) );
    zao21b U658 ( .A(INTDOORBELL), .B(DOORCNT_1), .C(n1618), .Y(DOORCNT1410_1)
         );
    zao21b U659 ( .A(INTDOORBELL), .B(DOORCNT_0), .C(n1619), .Y(DOORCNT1410_0)
         );
    zan2b U660 ( .A(n1667), .B(SWDBG), .Y(n1644) );
    zoa211b U661 ( .A(INTASYNC_S), .B(QHASYNCINT), .C(INTASYNC_EN), .D(n1645), 
        .Y(QHASYNCINT1448) );
    znd2b U662 ( .A(INTASYNC), .B(LTINT_PCLK), .Y(n1645) );
    zivb U663 ( .A(n1682), .Y(HEADSEEN_PRE) );
    zmux21lb U664 ( .A(HEADSEEN1), .B(HEADSEEN2), .S(CACHE_SEL_PRE), .Y(n1682)
         );
    zoai21b U665 ( .A(n1633), .B(n1634), .C(n1635), .Y(EHCISLEEP1231) );
    zan3b U666 ( .A(EHCIRESTART_SYNC), .B(ASYNCSM_0), .C(START_EVENT), .Y(
        n1633) );
    zmux21lb U667 ( .A(ASYNC_EMPTY1), .B(ASYNC_EMPTY2), .S(CACHE_SEL), .Y(
        n1635) );
    zor2b U668 ( .A(QCMDSTART1), .B(QCMDSTART2), .Y(TRANEXED1268) );
    zor2b U669 ( .A(EHCIRESTART), .B(EHCIRESTART_T), .Y(EHCIRESTART_SYNC313)
         );
    zxo2b U670 ( .A(QH_ACT2), .B(n1661), .Y(QH_ACT_SEL552) );
    zivb U671 ( .A(n1629), .Y(n1623) );
    zan2b U672 ( .A(n1819), .B(n1740), .Y(n1624) );
    zivb U673 ( .A(n1732), .Y(n1819) );
    zivb U674 ( .A(INTDOORBELL), .Y(n1740) );
    zao32b U675 ( .A(QHIDLE2), .B(n1774), .C(CACHEHIT2), .D(n1818), .E(
        CACHEHIT1), .Y(n1625) );
    zivb U676 ( .A(n1676), .Y(CACHEHIT2) );
    zivb U677 ( .A(n1674), .Y(CACHEHIT1) );
    zan3b U678 ( .A(n1636), .B(n1637), .C(n1638), .Y(EXE_HALT_pre) );
    znd2b U679 ( .A(RUN), .B(RUN_T), .Y(n1636) );
    zivb U680 ( .A(n1670), .Y(n1637) );
    zor2b U681 ( .A(n1640), .B(n1632), .Y(n1670) );
    zivb U682 ( .A(ASYNCSMNXT_1), .Y(n1638) );
    zoai211b U683 ( .A(PCIEND), .B(n1629), .C(n1630), .D(n1631), .Y(
        ASYNCSMNXT_1) );
    zivb U684 ( .A(n1636), .Y(RUN_ASYNC) );
    zoa211b U685 ( .A(n1652), .B(n1617), .C(n1648), .D(n1653), .Y(ASYNCSMNXT_4
        ) );
    zan2b U686 ( .A(n1672), .B(n1620), .Y(n1652) );
    zao32b U687 ( .A(n1648), .B(n1649), .C(n1650), .D(n1616), .E(n1651), .Y(
        ASYNCSMNXT_3) );
    zivb U688 ( .A(n1691), .Y(n1648) );
    zao21b U689 ( .A(EXE_HALT), .B(n1662), .C(GEN_PERR), .Y(n1691) );
    zivb U690 ( .A(SWDBG), .Y(n1662) );
    zor2b U691 ( .A(QHCIREQ1), .B(QHCIREQ2), .Y(n1649) );
    zao21b U692 ( .A(n1672), .B(n1620), .C(n1617), .Y(n1650) );
    zivb U693 ( .A(n1686), .Y(n1672) );
    zor2b U694 ( .A(PARSEQHEND2), .B(PARSEQHEND1), .Y(n1651) );
    zivb U695 ( .A(n1649), .Y(n1653) );
    zivb U696 ( .A(n1651), .Y(n1622) );
    zcx3b U697 ( .A(START_EVENT), .B(n1641), .C(n1642), .D(n1643), .Y(
        RECLAMATION1194) );
    zmux21lb U698 ( .A(QTDEXE1), .B(QTDEXE2), .S(QH_ACT2), .Y(n1642) );
    zao21b U699 ( .A(TRANEXED), .B(SWDBG), .C(GEN_PERR), .Y(RUN_C) );
    zao21b U700 ( .A(NAKCNTSM[0]), .B(n1656), .C(n1657), .Y(NAKCNTSMNXT[0]) );
    zivb U701 ( .A(n1779), .Y(HEADSEEN) );
    zan2b U702 ( .A(n1658), .B(NAKCNTSM[0]), .Y(NAKCNTSMNXT[1]) );
    zmux21lb U703 ( .A(n1779), .B(START_EVENT), .S(NAKCNTSM[1]), .Y(n1658) );
    zoai21b U704 ( .A(ASYNCSMNXT_0), .B(ASYNC_ACT), .C(n1621), .Y(START_EVENT)
         );
    zivb U705 ( .A(START_EVENT), .Y(n1656) );
    zivb U706 ( .A(ASYNCSMNXT_0), .Y(n1641) );
    zivb U707 ( .A(n1820), .Y(QH_CACHE_EN2) );
    zor2b U708 ( .A(n1689), .B(n1734), .Y(n1820) );
    zivb U709 ( .A(n1822), .Y(QH_CACHE_EN1) );
    zor2b U710 ( .A(CACHE_SEL), .B(n1689), .Y(n1822) );
    zan2b U711 ( .A(n1640), .B(QH_ACT2), .Y(ASYNC_EXE2) );
    zivb U712 ( .A(QHIDLE2), .Y(n1640) );
    zan2b U713 ( .A(n1632), .B(QH_ACT1), .Y(ASYNC_EXE1) );
    zivb U714 ( .A(QHIDLE1), .Y(n1632) );
    zor2b U715 ( .A(n1614), .B(QH_PARSE_GO2_T), .Y(QH_PARSE_GO2) );
    zor2b U716 ( .A(n1613), .B(QH_PARSE_GO1_T), .Y(QH_PARSE_GO1) );
    zivb U717 ( .A(PHASENXT_ParseQH), .Y(n1824) );
    zivb U718 ( .A(n1680), .Y(CACHE_SEL_PRE) );
    zivb U719 ( .A(PCIEND), .Y(n1639) );
    zivb U720 ( .A(QHCIREQ1), .Y(n1664) );
    zivb U721 ( .A(QHCIREQ2), .Y(n1665) );
    zdffrb NAKCNTSM_reg_1 ( .CK(PCICLK), .D(NAKCNTSMNXT[1]), .R(TRST_), .Q(
        NAKCNTSM[1]), .QN(n1666) );
    zdffqrb NAKCNTSM_reg_0 ( .CK(PCICLK), .D(NAKCNTSMNXT[0]), .R(TRST_), .Q(
        NAKCNTSM[0]) );
    zdffqrb CACHE_ADDR1_reg_26 ( .CK(PCICLK), .D(CACHE_ADDR1721_26), .R(TRST_), 
        .Q(CACHE_ADDR1[26]) );
    zdffqrb CACHE_ADDR1_reg_25 ( .CK(PCICLK), .D(CACHE_ADDR1721_25), .R(TRST_), 
        .Q(CACHE_ADDR1[25]) );
    zivb U722 ( .A(CACHE_ADDR1[25]), .Y(n1720) );
    zdffqrb CACHE_ADDR1_reg_24 ( .CK(PCICLK), .D(CACHE_ADDR1721_24), .R(TRST_), 
        .Q(CACHE_ADDR1[24]) );
    zivb U723 ( .A(CACHE_ADDR1[24]), .Y(n1722) );
    zdffqrb CACHE_ADDR1_reg_23 ( .CK(PCICLK), .D(CACHE_ADDR1721_23), .R(TRST_), 
        .Q(CACHE_ADDR1[23]) );
    zdffqrb CACHE_ADDR1_reg_22 ( .CK(PCICLK), .D(CACHE_ADDR1721_22), .R(TRST_), 
        .Q(CACHE_ADDR1[22]) );
    zdffqrb CACHE_ADDR1_reg_21 ( .CK(PCICLK), .D(CACHE_ADDR1721_21), .R(TRST_), 
        .Q(CACHE_ADDR1[21]) );
    zivb U724 ( .A(CACHE_ADDR1[21]), .Y(n1723) );
    zdffqrb CACHE_ADDR1_reg_20 ( .CK(PCICLK), .D(CACHE_ADDR1721_20), .R(TRST_), 
        .Q(CACHE_ADDR1[20]) );
    zivb U725 ( .A(CACHE_ADDR1[20]), .Y(n1715) );
    zdffqrb CACHE_ADDR1_reg_19 ( .CK(PCICLK), .D(CACHE_ADDR1721_19), .R(TRST_), 
        .Q(CACHE_ADDR1[19]) );
    zivb U726 ( .A(CACHE_ADDR1[19]), .Y(n1717) );
    zdffqrb CACHE_ADDR1_reg_18 ( .CK(PCICLK), .D(CACHE_ADDR1721_18), .R(TRST_), 
        .Q(CACHE_ADDR1[18]) );
    zdffqrb CACHE_ADDR1_reg_17 ( .CK(PCICLK), .D(CACHE_ADDR1721_17), .R(TRST_), 
        .Q(CACHE_ADDR1[17]) );
    zdffqrb CACHE_ADDR1_reg_16 ( .CK(PCICLK), .D(CACHE_ADDR1721_16), .R(TRST_), 
        .Q(CACHE_ADDR1[16]) );
    zdffqrb CACHE_ADDR1_reg_15 ( .CK(PCICLK), .D(CACHE_ADDR1721_15), .R(TRST_), 
        .Q(CACHE_ADDR1[15]) );
    zdffqrb CACHE_ADDR1_reg_14 ( .CK(PCICLK), .D(CACHE_ADDR1721_14), .R(TRST_), 
        .Q(CACHE_ADDR1[14]) );
    zdffqrb CACHE_ADDR1_reg_13 ( .CK(PCICLK), .D(CACHE_ADDR1721_13), .R(TRST_), 
        .Q(CACHE_ADDR1[13]) );
    zivb U727 ( .A(CACHE_ADDR1[13]), .Y(n1716) );
    zdffqrb CACHE_ADDR1_reg_12 ( .CK(PCICLK), .D(CACHE_ADDR1721_12), .R(TRST_), 
        .Q(CACHE_ADDR1[12]) );
    zivb U728 ( .A(CACHE_ADDR1[12]), .Y(n1721) );
    zdffqrb CACHE_ADDR1_reg_11 ( .CK(PCICLK), .D(CACHE_ADDR1721_11), .R(TRST_), 
        .Q(CACHE_ADDR1[11]) );
    zdffqrb CACHE_ADDR1_reg_10 ( .CK(PCICLK), .D(CACHE_ADDR1721_10), .R(TRST_), 
        .Q(CACHE_ADDR1[10]) );
    zdffqrb CACHE_ADDR1_reg_9 ( .CK(PCICLK), .D(CACHE_ADDR1721_9), .R(TRST_), 
        .Q(CACHE_ADDR1[9]) );
    zdffqrb CACHE_ADDR1_reg_8 ( .CK(PCICLK), .D(CACHE_ADDR1721_8), .R(TRST_), 
        .Q(CACHE_ADDR1[8]) );
    zivb U729 ( .A(CACHE_ADDR1[8]), .Y(n1713) );
    zdffqrb CACHE_ADDR1_reg_7 ( .CK(PCICLK), .D(CACHE_ADDR1721_7), .R(TRST_), 
        .Q(CACHE_ADDR1[7]) );
    zivb U730 ( .A(CACHE_ADDR1[7]), .Y(n1724) );
    zdffqrb CACHE_ADDR1_reg_6 ( .CK(PCICLK), .D(CACHE_ADDR1721_6), .R(TRST_), 
        .Q(CACHE_ADDR1[6]) );
    zivb U731 ( .A(CACHE_ADDR1[6]), .Y(n1718) );
    zdffqrb CACHE_ADDR1_reg_5 ( .CK(PCICLK), .D(CACHE_ADDR1721_5), .R(TRST_), 
        .Q(CACHE_ADDR1[5]) );
    zivb U732 ( .A(CACHE_ADDR1[5]), .Y(n1719) );
    zdffqrb CACHE_ADDR1_reg_4 ( .CK(PCICLK), .D(CACHE_ADDR1721_4), .R(TRST_), 
        .Q(CACHE_ADDR1[4]) );
    zdffqrb CACHE_ADDR1_reg_3 ( .CK(PCICLK), .D(CACHE_ADDR1721_3), .R(TRST_), 
        .Q(CACHE_ADDR1[3]) );
    zdffqrb CACHE_ADDR1_reg_2 ( .CK(PCICLK), .D(CACHE_ADDR1721_2), .R(TRST_), 
        .Q(CACHE_ADDR1[2]) );
    zivb U733 ( .A(CACHE_ADDR1[2]), .Y(n1725) );
    zdffqrb CACHE_ADDR1_reg_1 ( .CK(PCICLK), .D(CACHE_ADDR1721_1), .R(TRST_), 
        .Q(CACHE_ADDR1[1]) );
    zivb U734 ( .A(CACHE_ADDR1[1]), .Y(n1712) );
    zdffqrb CACHE_ADDR1_reg_0 ( .CK(PCICLK), .D(CACHE_ADDR1721_0), .R(TRST_), 
        .Q(CACHE_ADDR1[0]) );
    zivb U735 ( .A(CACHE_ADDR1[0]), .Y(n1714) );
    zdffqrb CACHE_ADDR2_reg_26 ( .CK(PCICLK), .D(CACHE_ADDR2759_26), .R(TRST_), 
        .Q(CACHE_ADDR2[26]) );
    zivb U736 ( .A(CACHE_ADDR2[26]), .Y(n1701) );
    zdffqrb CACHE_ADDR2_reg_25 ( .CK(PCICLK), .D(CACHE_ADDR2759_25), .R(TRST_), 
        .Q(CACHE_ADDR2[25]) );
    zdffqrb CACHE_ADDR2_reg_24 ( .CK(PCICLK), .D(CACHE_ADDR2759_24), .R(TRST_), 
        .Q(CACHE_ADDR2[24]) );
    zdffqrb CACHE_ADDR2_reg_23 ( .CK(PCICLK), .D(CACHE_ADDR2759_23), .R(TRST_), 
        .Q(CACHE_ADDR2[23]) );
    zdffqrb CACHE_ADDR2_reg_22 ( .CK(PCICLK), .D(CACHE_ADDR2759_22), .R(TRST_), 
        .Q(CACHE_ADDR2[22]) );
    zivb U737 ( .A(CACHE_ADDR2[22]), .Y(n1704) );
    zdffqrb CACHE_ADDR2_reg_21 ( .CK(PCICLK), .D(CACHE_ADDR2759_21), .R(TRST_), 
        .Q(CACHE_ADDR2[21]) );
    zivb U738 ( .A(CACHE_ADDR2[21]), .Y(n1692) );
    zdffqrb CACHE_ADDR2_reg_20 ( .CK(PCICLK), .D(CACHE_ADDR2759_20), .R(TRST_), 
        .Q(CACHE_ADDR2[20]) );
    zivb U739 ( .A(CACHE_ADDR2[20]), .Y(n1702) );
    zdffqrb CACHE_ADDR2_reg_19 ( .CK(PCICLK), .D(CACHE_ADDR2759_19), .R(TRST_), 
        .Q(CACHE_ADDR2[19]) );
    zivb U740 ( .A(CACHE_ADDR2[19]), .Y(n1695) );
    zdffqrb CACHE_ADDR2_reg_18 ( .CK(PCICLK), .D(CACHE_ADDR2759_18), .R(TRST_), 
        .Q(CACHE_ADDR2[18]) );
    zivb U741 ( .A(CACHE_ADDR2[18]), .Y(n1697) );
    zdffqrb CACHE_ADDR2_reg_17 ( .CK(PCICLK), .D(CACHE_ADDR2759_17), .R(TRST_), 
        .Q(CACHE_ADDR2[17]) );
    zivb U742 ( .A(CACHE_ADDR2[17]), .Y(n1699) );
    zdffqrb CACHE_ADDR2_reg_16 ( .CK(PCICLK), .D(CACHE_ADDR2759_16), .R(TRST_), 
        .Q(CACHE_ADDR2[16]) );
    zdffqrb CACHE_ADDR2_reg_15 ( .CK(PCICLK), .D(CACHE_ADDR2759_15), .R(TRST_), 
        .Q(CACHE_ADDR2[15]) );
    zivb U743 ( .A(CACHE_ADDR2[15]), .Y(n1705) );
    zdffqrb CACHE_ADDR2_reg_14 ( .CK(PCICLK), .D(CACHE_ADDR2759_14), .R(TRST_), 
        .Q(CACHE_ADDR2[14]) );
    zivb U744 ( .A(CACHE_ADDR2[14]), .Y(n1693) );
    zdffqrb CACHE_ADDR2_reg_13 ( .CK(PCICLK), .D(CACHE_ADDR2759_13), .R(TRST_), 
        .Q(CACHE_ADDR2[13]) );
    zivb U745 ( .A(CACHE_ADDR2[13]), .Y(n1694) );
    zdffqrb CACHE_ADDR2_reg_12 ( .CK(PCICLK), .D(CACHE_ADDR2759_12), .R(TRST_), 
        .Q(CACHE_ADDR2[12]) );
    zivb U746 ( .A(CACHE_ADDR2[12]), .Y(n1700) );
    zdffqrb CACHE_ADDR2_reg_11 ( .CK(PCICLK), .D(CACHE_ADDR2759_11), .R(TRST_), 
        .Q(CACHE_ADDR2[11]) );
    zdffqrb CACHE_ADDR2_reg_10 ( .CK(PCICLK), .D(CACHE_ADDR2759_10), .R(TRST_), 
        .Q(CACHE_ADDR2[10]) );
    zdffqrb CACHE_ADDR2_reg_9 ( .CK(PCICLK), .D(CACHE_ADDR2759_9), .R(TRST_), 
        .Q(CACHE_ADDR2[9]) );
    zdffqrb CACHE_ADDR2_reg_8 ( .CK(PCICLK), .D(CACHE_ADDR2759_8), .R(TRST_), 
        .Q(CACHE_ADDR2[8]) );
    zdffqrb CACHE_ADDR2_reg_7 ( .CK(PCICLK), .D(CACHE_ADDR2759_7), .R(TRST_), 
        .Q(CACHE_ADDR2[7]) );
    zdffqrb CACHE_ADDR2_reg_6 ( .CK(PCICLK), .D(CACHE_ADDR2759_6), .R(TRST_), 
        .Q(CACHE_ADDR2[6]) );
    zdffqrb CACHE_ADDR2_reg_5 ( .CK(PCICLK), .D(CACHE_ADDR2759_5), .R(TRST_), 
        .Q(CACHE_ADDR2[5]) );
    zdffqrb CACHE_ADDR2_reg_4 ( .CK(PCICLK), .D(CACHE_ADDR2759_4), .R(TRST_), 
        .Q(CACHE_ADDR2[4]) );
    zivb U747 ( .A(CACHE_ADDR2[4]), .Y(n1703) );
    zdffqrb CACHE_ADDR2_reg_3 ( .CK(PCICLK), .D(CACHE_ADDR2759_3), .R(TRST_), 
        .Q(CACHE_ADDR2[3]) );
    zivb U748 ( .A(CACHE_ADDR2[3]), .Y(n1698) );
    zdffqrb CACHE_ADDR2_reg_2 ( .CK(PCICLK), .D(CACHE_ADDR2759_2), .R(TRST_), 
        .Q(CACHE_ADDR2[2]) );
    zivb U749 ( .A(CACHE_ADDR2[2]), .Y(n1696) );
    zdffqrb CACHE_ADDR2_reg_1 ( .CK(PCICLK), .D(CACHE_ADDR2759_1), .R(TRST_), 
        .Q(CACHE_ADDR2[1]) );
    zdffqrb CACHE_ADDR2_reg_0 ( .CK(PCICLK), .D(CACHE_ADDR2759_0), .R(TRST_), 
        .Q(CACHE_ADDR2[0]) );
    zdffqrb DOORCNT_reg_1 ( .CK(PCICLK), .D(DOORCNT1410_1), .R(TRST_), .Q(
        DOORCNT_1) );
    zivb U750 ( .A(DOORCNT_1), .Y(n1738) );
    zdffqrb DOORCNT_reg_0 ( .CK(PCICLK), .D(DOORCNT1410_0), .R(TRST_), .Q(
        DOORCNT_0) );
    zivb U751 ( .A(DOORCNT_0), .Y(n1737) );
    zdffqsb FROZEN_reg ( .CK(PCICLK), .D(FROZEN1366), .S(TRST_), .Q(FROZEN) );
    zdffqrb ASYNCSM_reg_1 ( .CK(PCICLK), .D(ASYNCSMNXT_1), .R(TRST_), .Q(
        ASYNCSM_1) );
    zivb U752 ( .A(ASYNCSM_1), .Y(n1688) );
    zdffqrb EHCIRESTART_T_reg ( .CK(PCICLK), .D(EHCIRESTART), .R(TRST_), .Q(
        EHCIRESTART_T) );
    zdffqrb QHASYNCINT_reg ( .CK(PCICLK), .D(QHASYNCINT1448), .R(TRST_), .Q(
        QHASYNCINT) );
    zdffqrb QH_PARSE_GO1_T_reg ( .CK(PCICLK), .D(n1613), .R(TRST_), .Q(
        QH_PARSE_GO1_T) );
    zdffqrb HEADSEEN_T_reg ( .CK(PCICLK), .D(HEADSEEN_PRE), .R(TRST_), .Q(
        HEADSEEN_T) );
    zdffqrb EHCISLEEP_reg ( .CK(PCICLK), .D(EHCISLEEP1231), .R(TRST_), .Q(
        EHCISLEEP) );
    zivb U753 ( .A(EHCISLEEP), .Y(n1634) );
    zdffsb ASYNCSM_reg_0 ( .CK(PCICLK), .D(ASYNCSMNXT_0), .S(TRST_), .Q(
        ASYNCSM_0), .QN(ASYNC_ACT) );
    zdffqrb TRANEXED_reg ( .CK(PCICLK), .D(TRANEXED1268), .R(TRST_), .Q(
        TRANEXED) );
    zdffqrb EHCIRESTART_SYNC_reg ( .CK(PCICLK), .D(EHCIRESTART_SYNC313), .R(
        TRST_), .Q(EHCIRESTART_SYNC) );
    zivb U754 ( .A(EHCIRESTART_SYNC), .Y(n1739) );
    zdffrb QH_ACT_SEL_reg ( .CK(PCICLK), .D(QH_ACT_SEL552), .R(TRST_), .Q(
        QH_ACT2), .QN(QH_ACT1) );
    zdffqrb ASYNCSM_reg_2 ( .CK(PCICLK), .D(PHASENXT_ParseQH), .R(TRST_), .Q(
        PHASE_ParseQH) );
    zivb U755 ( .A(PHASE_ParseQH), .Y(n1689) );
    zdffqrb CACHE_SEL_reg ( .CK(PCICLK), .D(CACHE_SEL_PRE), .R(TRST_), .Q(
        CACHE_SEL) );
    zivb U756 ( .A(CACHE_SEL), .Y(n1734) );
    zdffqrb RUN_T_reg ( .CK(PCICLK), .D(RUN), .R(TRST_), .Q(RUN_T) );
    zdffqsb EXE_HALT_reg ( .CK(PCICLK), .D(EXE_HALT_pre), .S(TRST_), .Q(
        EXE_HALT) );
    zdffqrb ASYNCSM_reg_4 ( .CK(PCICLK), .D(ASYNCSMNXT_4), .R(TRST_), .Q(
        ASYNCSM_4) );
    zivb U757 ( .A(ASYNCSM_4), .Y(n1685) );
    zdffqrb HEADSEEN_2T_reg ( .CK(PCICLK), .D(HEADSEEN), .R(TRST_), .Q(
        HEADSEEN_2T) );
    zdffqrb ASYNCSM_reg_3 ( .CK(PCICLK), .D(ASYNCSMNXT_3), .R(TRST_), .Q(
        ASYNCSM_3) );
    zivb U758 ( .A(ASYNCSM_3), .Y(n1687) );
    zdffqrb RECLAMATION_reg ( .CK(PCICLK), .D(RECLAMATION1194), .R(TRST_), .Q(
        RECLAMATION) );
    zdffqrb QH_PARSE_GO2_T_reg ( .CK(PCICLK), .D(n1614), .R(TRST_), .Q(
        QH_PARSE_GO2_T) );
    zdffqrb LIST_SEL_T_reg ( .CK(PCICLK), .D(LIST_SEL), .R(TRST_), .Q(
        LIST_SEL_T) );
    zaoi21b U759 ( .A(n1820), .B(n1821), .C(n1665), .Y(QHCIGNT2) );
    zaoi21b U760 ( .A(n1822), .B(n1823), .C(n1664), .Y(QHCIGNT1) );
    znr3b U761 ( .A(PHASE_ParseQH), .B(n1824), .C(CACHE_SEL_PRE), .Y(n1613) );
    znr3b U762 ( .A(PHASE_ParseQH), .B(n1824), .C(n1680), .Y(n1614) );
    znr2b U763 ( .A(n1737), .B(n1738), .Y(INTASYNC_S) );
    znr3b U764 ( .A(ASYNCSM_1), .B(n1689), .C(n1733), .Y(n1616) );
    znr3b U765 ( .A(ASYNCSM_1), .B(n1687), .C(n1690), .Y(n1617) );
    znr2b U766 ( .A(n1640), .B(n1740), .Y(n1618) );
    znr2b U767 ( .A(n1632), .B(n1740), .Y(n1619) );
    zmux21hb U768 ( .A(n1671), .B(n1670), .S(EHCISLEEP), .Y(n1620) );
    zao222b U769 ( .A(n1616), .B(n1622), .C(PCIEND), .D(n1623), .E(n1624), .F(
        n1625), .Y(PHASENXT_ParseQH) );
    zor3b U770 ( .A(n1626), .B(n1627), .C(n1628), .Y(ASYNCSMNXT_0) );
    zao211b U771 ( .A(ASYNCSM_1), .B(n1639), .C(QHCIGNT1), .D(QHCIGNT2), .Y(
        EHCIREQ) );
    zoa21d U772 ( .A(n1644), .B(FROZEN), .C(n1636), .Y(FROZEN1366) );
    zoa21d U773 ( .A(EHCISLEEP), .B(n1659), .C(n1660), .Y(n1628) );
    zoa21d U774 ( .A(RUN), .B(n1662), .C(n1663), .Y(n1661) );
    zoa21d U775 ( .A(NAKCNTSM[0]), .B(HEADSEEN), .C(n1666), .Y(n1657) );
    zoa21d U776 ( .A(CACHEHIT2), .B(n1669), .C(QHIDLE2), .Y(n1668) );
    zor3b U777 ( .A(ASYNC_ACT), .B(n1678), .C(n1683), .Y(n1684) );
    zor4b U778 ( .A(ASYNCSM_0), .B(PHASE_ParseQH), .C(n1685), .D(n1678), .Y(
        n1686) );
    zor6b U779 ( .A(n1706), .B(n1707), .C(n1708), .D(n1709), .E(n1710), .F(
        n1711), .Y(n1676) );
    zor6b U780 ( .A(n1726), .B(n1727), .C(n1728), .D(n1729), .E(n1730), .F(
        n1731), .Y(n1674) );
    zor4b U781 ( .A(EHCISLEEP), .B(n1686), .C(n1691), .D(n1636), .Y(n1732) );
    zor4b U782 ( .A(ASYNCSM_3), .B(ASYNCSM_4), .C(ASYNCSM_0), .D(n1691), .Y(
        n1733) );
    zor3b U783 ( .A(PHASE_ParseQH), .B(n1688), .C(n1733), .Y(n1629) );
    zor3b U784 ( .A(ASYNCSM_0), .B(CACHE_INVALID2), .C(n1618), .Y(n1742) );
    zor3b U785 ( .A(ASYNCSM_0), .B(CACHE_INVALID1), .C(n1619), .Y(n1748) );
    zcx8d U786 ( .A(ASYNC_EN), .B(n1670), .C(n1780), .D(n1781), .E(n1782), .Y(
        n1671) );
    zao222b U787 ( .A(ASYNCSM_1), .B(ASYNCSM_3), .C(n1683), .D(ASYNCSM_0), .E(
        n1784), .F(n1636), .Y(n1626) );
    zao211b U788 ( .A(PHASE_ParseQH), .B(ASYNCSM_4), .C(n1677), .D(n1691), .Y(
        n1627) );
    zan4b U789 ( .A(n1787), .B(n1788), .C(n1789), .D(n1790), .Y(n1786) );
    zan4b U790 ( .A(n1792), .B(n1793), .C(n1794), .D(n1795), .Y(n1791) );
    zor4b U791 ( .A(n1755), .B(n1756), .C(n1753), .D(n1754), .Y(n1709) );
    zor6b U792 ( .A(n1760), .B(n1761), .C(n1762), .D(n1757), .E(n1758), .F(
        n1759), .Y(n1710) );
    zan4b U793 ( .A(n1803), .B(n1804), .C(n1805), .D(n1806), .Y(n1802) );
    zan4b U794 ( .A(n1808), .B(n1809), .C(n1810), .D(n1811), .Y(n1807) );
    zor4b U795 ( .A(n1765), .B(n1766), .C(n1763), .D(n1764), .Y(n1729) );
    zor6b U796 ( .A(n1770), .B(n1771), .C(n1772), .D(n1767), .E(n1768), .F(
        n1769), .Y(n1730) );
    zoa21d U797 ( .A(ASYNC_EN), .B(n1640), .C(QHIDLE1), .Y(n1818) );
    zoa21d U798 ( .A(n1669), .B(n1740), .C(RUN_ASYNC), .Y(n1780) );
    zind2d U799 ( .A(LIST_SEL_T), .B(LIST_SEL), .Y(n1621) );
    zind2d U800 ( .A(HEADSEEN_2T), .B(RECLAMATION), .Y(n1643) );
    zor3b U801 ( .A(EHCISLEEP), .B(n1659), .C(n1636), .Y(n1825) );
    zor3b U802 ( .A(n1773), .B(n1732), .C(CACHE_HIT), .Y(n1631) );
    zao211b U803 ( .A(n1739), .B(n1825), .C(n1691), .D(n1684), .Y(n1630) );
    zao211b U804 ( .A(n1638), .B(n1824), .C(n1775), .D(n1685), .Y(n1681) );
    zor3b U805 ( .A(PHASE_ParseQH), .B(n1687), .C(n1783), .Y(n1821) );
    zor3b U806 ( .A(PHASE_ParseQH), .B(n1687), .C(n1826), .Y(n1823) );
    zor3b U807 ( .A(QHIDLE2), .B(CACHEHIT1), .C(n1669), .Y(n1781) );
endmodule


module HS_PCICTL ( LDW, PCI1WAIT, HCIMRDY, RDYACK, HCICOMPL, PCIEND, MABORTS, 
    TABORTR, GEN_PERR, HCIGNT, PCICLK, TRST_, PAROPT, PERRS, SERRS, PMSTR, 
    MADDR, EDWNUM, DWCNT, HCIMWR, EDWOFFSET, UGNTI_, ATPG_ENI );
output [15:0] LDW;
input  [3:0] EDWNUM;
output [3:0] DWCNT;
input  [3:0] EDWOFFSET;
input  PCI1WAIT, RDYACK, MABORTS, TABORTR, HCIGNT, PCICLK, TRST_, PAROPT, 
    PERRS, SERRS, PMSTR, HCIMWR, UGNTI_, ATPG_ENI;
output HCIMRDY, HCICOMPL, PCIEND, GEN_PERR, MADDR;
    wire PCISMNXT_2, SPAREO6, LDW597_12, LDW597_1, LDW597_8, SPAREO0_, SPAREO8, 
        PCIEND635, LDW597_15, LDW597_6, DWCNT513_0, DWCNT497_1, DWCNT_N_1, 
        SPAREO1, SPAREO9, PCIEND_RST_, DWCNT497_0, DWCNT_N_0, SPAREO0, 
        DWCNT513_1, PCISMNXT_3, LDW597_14, LDW597_7, LDW597_13, LDW597_0, 
        SPAREO7, LDW597_9, PCISMNXT_1, SPAREO5, LDW597_11, LDW597_2, PCISM_0, 
        LDW597_5, DWCNT513_3, DWCNT_N_2, SPAREO2, DWCNT497_2, DWINC, MADDR555, 
        DWCNT_N_3, SPAREO3, SPAREO1_, DWCNT497_3, PCISM_1, PCISMNXT_0, 
        DWCNT513_2, LDW597_4, LDW597_10, LDW597_3, SPAREO4, n736, n737, n738, 
        n739, n740, n741, n742, n743, n744, n745, n746, add_105_carry_2, 
        add_105_carry_3, n747, n748, n749, n750, n751, n752, n753, n754, n755, 
        n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, 
        n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
        n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, 
        n792, n793, n794, n795, n796, n797, n798, n799;
    zdffrb SPARE550 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE559 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb SPARE557 ( .A(SPAREO4), .Y(SPAREO5) );
    zdffrb SPARE551 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    znr3b SPARE556 ( .A(SPAREO2), .B(DWINC), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE558 ( .A(SPAREO5), .Y(SPAREO6) );
    zaoi211b SPARE553 ( .A(SPAREO4), .B(PCIEND_RST_), .C(SPAREO6), .D(1'b0), 
        .Y(SPAREO8) );
    zoai21b SPARE554 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zoai21b SPARE555 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE552 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    znd2b U229 ( .A(EDWOFFSET[1]), .B(n747), .Y(n751) );
    znd2b U230 ( .A(n753), .B(n754), .Y(n747) );
    znd2b U231 ( .A(DWCNT[1]), .B(n750), .Y(n752) );
    znr2b U232 ( .A(n761), .B(n758), .Y(n757) );
    zaoi21b U233 ( .A(n746), .B(n760), .C(n759), .Y(n761) );
    znr2b U234 ( .A(n746), .B(n760), .Y(n758) );
    zxo2b U235 ( .A(n748), .B(EDWOFFSET[3]), .Y(n756) );
    zor2b U236 ( .A(n787), .B(n778), .Y(n794) );
    zor2b U237 ( .A(n786), .B(n788), .Y(n789) );
    zxo2b U238 ( .A(n750), .B(n749), .Y(DWCNT_N_1) );
    zivb U239 ( .A(n754), .Y(n750) );
    znd2b U240 ( .A(EDWOFFSET[0]), .B(DWCNT[0]), .Y(n754) );
    zxo2b U241 ( .A(EDWOFFSET[1]), .B(DWCNT[1]), .Y(n749) );
    zxo2b U242 ( .A(n755), .B(n746), .Y(DWCNT_N_2) );
    zxo2b U243 ( .A(n759), .B(DWCNT[2]), .Y(n755) );
    zivb U244 ( .A(EDWOFFSET[2]), .Y(n759) );
    zor2b U245 ( .A(DWCNT_N_3), .B(n786), .Y(n793) );
    zxo2b U246 ( .A(n756), .B(n757), .Y(DWCNT_N_3) );
    zivb U247 ( .A(DWCNT_N_3), .Y(n788) );
    zxo2b U248 ( .A(EDWOFFSET[0]), .B(DWCNT[0]), .Y(DWCNT_N_0) );
    zmux21lb U249 ( .A(n785), .B(n795), .S(HCIMRDY), .Y(n799) );
    zor2b U250 ( .A(PCISM_1), .B(n796), .Y(n795) );
    zor2b U251 ( .A(PCISM_1), .B(HCIMRDY), .Y(n774) );
    zxo2b U252 ( .A(n775), .B(n787), .Y(n798) );
    zivb U253 ( .A(n774), .Y(n787) );
    znd2b U254 ( .A(PMSTR), .B(RDYACK), .Y(n778) );
    zivb U255 ( .A(n778), .Y(n796) );
    zoa211b U256 ( .A(PERRS), .B(SERRS), .C(PAROPT), .D(n767), .Y(n769) );
    zxo2b U257 ( .A(EDWNUM[0]), .B(DWCNT[0]), .Y(n784) );
    zxo2b U258 ( .A(EDWNUM[1]), .B(DWCNT[1]), .Y(n783) );
    zxo2b U259 ( .A(EDWNUM[3]), .B(DWCNT[3]), .Y(n782) );
    zxo2b U260 ( .A(EDWNUM[2]), .B(DWCNT[2]), .Y(n781) );
    zao22b U261 ( .A(DWCNT497_3), .B(n736), .C(n737), .D(DWCNT[3]), .Y(
        DWCNT513_3) );
    zxo2b U262 ( .A(add_105_carry_3), .B(DWCNT[3]), .Y(DWCNT497_3) );
    zao22b U263 ( .A(DWCNT497_2), .B(n736), .C(n737), .D(DWCNT[2]), .Y(
        DWCNT513_2) );
    zhadrb add_105_U1_1_2 ( .A(DWCNT[2]), .B(add_105_carry_2), .CO(
        add_105_carry_3), .S(DWCNT497_2) );
    zao22b U264 ( .A(DWCNT497_1), .B(n736), .C(n737), .D(DWCNT[1]), .Y(
        DWCNT513_1) );
    zhadrb add_105_U1_1_1 ( .A(DWCNT[1]), .B(DWCNT[0]), .CO(add_105_carry_2), 
        .S(DWCNT497_1) );
    zao22b U265 ( .A(DWCNT497_0), .B(n736), .C(n737), .D(DWCNT[0]), .Y(
        DWCNT513_0) );
    zivb U266 ( .A(n794), .Y(DWINC) );
    zan2b U267 ( .A(n738), .B(n742), .Y(LDW597_15) );
    zan2b U268 ( .A(n738), .B(n744), .Y(LDW597_14) );
    zan2b U269 ( .A(n739), .B(n742), .Y(LDW597_13) );
    zan2b U270 ( .A(n739), .B(n744), .Y(LDW597_12) );
    zan2b U271 ( .A(n740), .B(n742), .Y(LDW597_11) );
    zan2b U272 ( .A(n740), .B(n744), .Y(LDW597_10) );
    zan2b U273 ( .A(n741), .B(n742), .Y(LDW597_9) );
    zan2b U274 ( .A(n744), .B(n741), .Y(LDW597_8) );
    zan2b U275 ( .A(n738), .B(n743), .Y(LDW597_7) );
    zan2b U276 ( .A(n745), .B(n738), .Y(LDW597_6) );
    zan2b U277 ( .A(n739), .B(n743), .Y(LDW597_5) );
    zan2b U278 ( .A(n739), .B(n745), .Y(LDW597_4) );
    zivb U279 ( .A(DWCNT_N_2), .Y(n792) );
    zan2b U280 ( .A(n740), .B(n743), .Y(LDW597_3) );
    zan2b U281 ( .A(n740), .B(n745), .Y(LDW597_2) );
    zivb U282 ( .A(DWCNT_N_1), .Y(n791) );
    zan2b U283 ( .A(n743), .B(n741), .Y(LDW597_1) );
    zivb U284 ( .A(DWCNT_N_0), .Y(n790) );
    zan2b U285 ( .A(n745), .B(n741), .Y(LDW597_0) );
    zor2b U286 ( .A(HCIGNT), .B(ATPG_ENI), .Y(PCIEND_RST_) );
    zan2b U287 ( .A(PCISMNXT_0), .B(n767), .Y(PCIEND635) );
    zan2b U288 ( .A(n762), .B(n764), .Y(PCISMNXT_2) );
    zao32b U289 ( .A(n775), .B(n797), .C(n799), .D(n763), .E(n780), .Y(n764)
         );
    zivb U290 ( .A(PCI1WAIT), .Y(n780) );
    zan3b U291 ( .A(n762), .B(PCI1WAIT), .C(n763), .Y(PCISMNXT_1) );
    znr2b U292 ( .A(UGNTI_), .B(n767), .Y(MADDR555) );
    zoa211b U293 ( .A(n770), .B(n771), .C(n772), .D(n773), .Y(n765) );
    zor2b U294 ( .A(PCISMNXT_3), .B(n776), .Y(n766) );
    zivb U295 ( .A(HCIGNT), .Y(n776) );
    zivb U296 ( .A(n766), .Y(n762) );
    zao21b U297 ( .A(n768), .B(HCIMRDY), .C(GEN_PERR), .Y(HCICOMPL) );
    zivb U298 ( .A(n771), .Y(n768) );
    zdffqrb DWCNT_reg_3 ( .CK(PCICLK), .D(DWCNT513_3), .R(TRST_), .Q(DWCNT[3])
         );
    zivb U299 ( .A(DWCNT[3]), .Y(n748) );
    zdffqrb DWCNT_reg_2 ( .CK(PCICLK), .D(DWCNT513_2), .R(TRST_), .Q(DWCNT[2])
         );
    zivb U300 ( .A(DWCNT[2]), .Y(n760) );
    zdffqrb DWCNT_reg_1 ( .CK(PCICLK), .D(DWCNT513_1), .R(TRST_), .Q(DWCNT[1])
         );
    zivb U301 ( .A(DWCNT[1]), .Y(n753) );
    zdffqrb DWCNT_reg_0 ( .CK(PCICLK), .D(DWCNT513_0), .R(TRST_), .Q(DWCNT[0])
         );
    zivb U302 ( .A(DWCNT[0]), .Y(DWCNT497_0) );
    zdffqrb LDW_reg_15 ( .CK(PCICLK), .D(LDW597_15), .R(TRST_), .Q(LDW[15]) );
    zdffqrb LDW_reg_14 ( .CK(PCICLK), .D(LDW597_14), .R(TRST_), .Q(LDW[14]) );
    zdffqrb LDW_reg_13 ( .CK(PCICLK), .D(LDW597_13), .R(TRST_), .Q(LDW[13]) );
    zdffqrb LDW_reg_12 ( .CK(PCICLK), .D(LDW597_12), .R(TRST_), .Q(LDW[12]) );
    zdffqrb LDW_reg_11 ( .CK(PCICLK), .D(LDW597_11), .R(TRST_), .Q(LDW[11]) );
    zdffqrb LDW_reg_10 ( .CK(PCICLK), .D(LDW597_10), .R(TRST_), .Q(LDW[10]) );
    zdffqrb LDW_reg_9 ( .CK(PCICLK), .D(LDW597_9), .R(TRST_), .Q(LDW[9]) );
    zdffqrb LDW_reg_8 ( .CK(PCICLK), .D(LDW597_8), .R(TRST_), .Q(LDW[8]) );
    zdffqrb LDW_reg_7 ( .CK(PCICLK), .D(LDW597_7), .R(TRST_), .Q(LDW[7]) );
    zdffqrb LDW_reg_6 ( .CK(PCICLK), .D(LDW597_6), .R(TRST_), .Q(LDW[6]) );
    zdffqrb LDW_reg_5 ( .CK(PCICLK), .D(LDW597_5), .R(TRST_), .Q(LDW[5]) );
    zdffqrb LDW_reg_4 ( .CK(PCICLK), .D(LDW597_4), .R(TRST_), .Q(LDW[4]) );
    zdffqrb LDW_reg_3 ( .CK(PCICLK), .D(LDW597_3), .R(TRST_), .Q(LDW[3]) );
    zdffqrb LDW_reg_2 ( .CK(PCICLK), .D(LDW597_2), .R(TRST_), .Q(LDW[2]) );
    zdffqrb LDW_reg_1 ( .CK(PCICLK), .D(LDW597_1), .R(TRST_), .Q(LDW[1]) );
    zdffqrb LDW_reg_0 ( .CK(PCICLK), .D(LDW597_0), .R(TRST_), .Q(LDW[0]) );
    zdffqrb PCIEND_reg ( .CK(PCICLK), .D(PCIEND635), .R(PCIEND_RST_), .Q(
        PCIEND) );
    zdffqrb PCISM_reg_2 ( .CK(PCICLK), .D(PCISMNXT_2), .R(TRST_), .Q(HCIMRDY)
         );
    zivb U303 ( .A(HCIMRDY), .Y(n777) );
    zdffqrb PCISM_reg_3 ( .CK(PCICLK), .D(PCISMNXT_3), .R(TRST_), .Q(GEN_PERR)
         );
    zivb U304 ( .A(GEN_PERR), .Y(n797) );
    zdffqrb PCISM_reg_1 ( .CK(PCICLK), .D(PCISMNXT_1), .R(TRST_), .Q(PCISM_1)
         );
    zivb U305 ( .A(PCISM_1), .Y(n785) );
    zdffrb MADDR_reg ( .CK(PCICLK), .D(MADDR555), .R(TRST_), .Q(MADDR), .QN(
        n779) );
    zdffsb PCISM_reg_0 ( .CK(PCICLK), .D(PCISMNXT_0), .S(TRST_), .Q(PCISM_0), 
        .QN(n775) );
    znr2b U306 ( .A(PCISM_0), .B(n794), .Y(n736) );
    znr2b U307 ( .A(DWINC), .B(PCISM_0), .Y(n737) );
    znr2b U308 ( .A(n791), .B(n792), .Y(n738) );
    znr2b U309 ( .A(DWCNT_N_1), .B(n792), .Y(n739) );
    znr2b U310 ( .A(DWCNT_N_2), .B(n791), .Y(n740) );
    znr2b U311 ( .A(DWCNT_N_2), .B(DWCNT_N_1), .Y(n741) );
    znr2b U312 ( .A(n789), .B(n790), .Y(n742) );
    znr2b U313 ( .A(n790), .B(n793), .Y(n743) );
    znr2b U314 ( .A(DWCNT_N_0), .B(n789), .Y(n744) );
    znr2b U315 ( .A(DWCNT_N_0), .B(n793), .Y(n745) );
    zan2b U316 ( .A(n752), .B(n751), .Y(n746) );
    zoai22d U317 ( .A(HCIGNT), .B(PCISMNXT_3), .C(n765), .D(n766), .Y(
        PCISMNXT_0) );
    zor3b U318 ( .A(TABORTR), .B(MABORTS), .C(n769), .Y(PCISMNXT_3) );
    zor5b U319 ( .A(GEN_PERR), .B(PCISM_1), .C(PCISM_0), .D(n777), .E(n778), 
        .Y(n770) );
    zor3b U320 ( .A(GEN_PERR), .B(n775), .C(n774), .Y(n767) );
    zor4b U321 ( .A(n781), .B(n782), .C(n783), .D(n784), .Y(n771) );
    zor3b U322 ( .A(HCIMWR), .B(n787), .C(n778), .Y(n786) );
    zoa21d U323 ( .A(MADDR), .B(n767), .C(n797), .Y(n772) );
    zoa21d U324 ( .A(n777), .B(n785), .C(n798), .Y(n773) );
    zoai22d U325 ( .A(n767), .B(n779), .C(n768), .D(n770), .Y(n763) );
endmodule


module PHCI_CACHE ( LDW, ADI, PCICLK, TRST_, CACHE_EN, DW0, DW1, ATPG_ENI );
input  [15:0] LDW;
output [31:0] DW0;
input  [31:0] ADI;
output [31:0] DW1;
input  PCICLK, TRST_, CACHE_EN, ATPG_ENI;
    wire FLOPS_CLK_14, n_19, FLOPS_CLK_15, n_20, DNT_DW1_n126, DNT_DW1_n127, 
        DNT_DW0_n126, DNT_DW0_n127;
    zan2b U12 ( .A(CACHE_EN), .B(LDW[0]), .Y(n_20) );
    zan2b U13 ( .A(LDW[1]), .B(CACHE_EN), .Y(n_19) );
    zmux21hd U14 ( .A(n_19), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_15) );
    zmux21hd U15 ( .A(n_20), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_14) );
    zdffqrb DNT_DW1_Q_reg_31 ( .CK(DNT_DW1_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW1[31]) );
    zdffqrb DNT_DW1_Q_reg_30 ( .CK(DNT_DW1_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW1[30]) );
    zdffqrb DNT_DW1_Q_reg_29 ( .CK(DNT_DW1_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW1[29]) );
    zdffqrb DNT_DW1_Q_reg_28 ( .CK(DNT_DW1_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW1[28]) );
    zdffqrb DNT_DW1_Q_reg_27 ( .CK(DNT_DW1_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW1[27]) );
    zdffqrb DNT_DW1_Q_reg_26 ( .CK(DNT_DW1_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW1[26]) );
    zdffqrb DNT_DW1_Q_reg_25 ( .CK(DNT_DW1_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW1[25]) );
    zdffqrb DNT_DW1_Q_reg_24 ( .CK(DNT_DW1_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW1[24]) );
    zdffqrb DNT_DW1_Q_reg_23 ( .CK(DNT_DW1_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW1[23]) );
    zdffqrb DNT_DW1_Q_reg_22 ( .CK(DNT_DW1_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW1[22]) );
    zdffqrb DNT_DW1_Q_reg_21 ( .CK(DNT_DW1_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW1[21]) );
    zdffqrb DNT_DW1_Q_reg_20 ( .CK(DNT_DW1_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW1[20]) );
    zdffqrb DNT_DW1_Q_reg_19 ( .CK(DNT_DW1_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW1[19]) );
    zdffqrb DNT_DW1_Q_reg_18 ( .CK(DNT_DW1_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW1[18]) );
    zdffqrb DNT_DW1_Q_reg_17 ( .CK(DNT_DW1_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW1[17]) );
    zdffqrb DNT_DW1_Q_reg_16 ( .CK(DNT_DW1_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW1[16]) );
    zdffqrb DNT_DW1_Q_reg_15 ( .CK(DNT_DW1_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW1[15]) );
    zdffqrb DNT_DW1_Q_reg_14 ( .CK(DNT_DW1_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW1[14]) );
    zdffqrb DNT_DW1_Q_reg_13 ( .CK(DNT_DW1_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW1[13]) );
    zdffqrb DNT_DW1_Q_reg_12 ( .CK(DNT_DW1_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW1[12]) );
    zdffqrb DNT_DW1_Q_reg_11 ( .CK(DNT_DW1_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW1[11]) );
    zdffqrb DNT_DW1_Q_reg_10 ( .CK(DNT_DW1_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW1[10]) );
    zdffqrb DNT_DW1_Q_reg_9 ( .CK(DNT_DW1_n126), .D(ADI[9]), .R(TRST_), .Q(DW1
        [9]) );
    zdffqrb DNT_DW1_Q_reg_8 ( .CK(DNT_DW1_n126), .D(ADI[8]), .R(TRST_), .Q(DW1
        [8]) );
    zdffqrb DNT_DW1_Q_reg_7 ( .CK(DNT_DW1_n126), .D(ADI[7]), .R(TRST_), .Q(DW1
        [7]) );
    zdffqrb DNT_DW1_Q_reg_6 ( .CK(DNT_DW1_n126), .D(ADI[6]), .R(TRST_), .Q(DW1
        [6]) );
    zdffqrb DNT_DW1_Q_reg_5 ( .CK(DNT_DW1_n126), .D(ADI[5]), .R(TRST_), .Q(DW1
        [5]) );
    zdffqrb DNT_DW1_Q_reg_4 ( .CK(DNT_DW1_n126), .D(ADI[4]), .R(TRST_), .Q(DW1
        [4]) );
    zdffqrb DNT_DW1_Q_reg_3 ( .CK(DNT_DW1_n126), .D(ADI[3]), .R(TRST_), .Q(DW1
        [3]) );
    zdffqrb DNT_DW1_Q_reg_2 ( .CK(DNT_DW1_n126), .D(ADI[2]), .R(TRST_), .Q(DW1
        [2]) );
    zdffqrb DNT_DW1_Q_reg_1 ( .CK(DNT_DW1_n126), .D(ADI[1]), .R(TRST_), .Q(DW1
        [1]) );
    zdffqrb DNT_DW1_Q_reg_0 ( .CK(DNT_DW1_n126), .D(ADI[0]), .R(TRST_), .Q(DW1
        [0]) );
    zbfb DNT_DW1_U80 ( .A(FLOPS_CLK_15), .Y(DNT_DW1_n126) );
    zbfb DNT_DW1_U81 ( .A(FLOPS_CLK_15), .Y(DNT_DW1_n127) );
    zdffqrb DNT_DW0_Q_reg_31 ( .CK(DNT_DW0_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW0[31]) );
    zdffqrb DNT_DW0_Q_reg_30 ( .CK(DNT_DW0_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW0[30]) );
    zdffqrb DNT_DW0_Q_reg_29 ( .CK(DNT_DW0_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW0[29]) );
    zdffqrb DNT_DW0_Q_reg_28 ( .CK(DNT_DW0_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW0[28]) );
    zdffqrb DNT_DW0_Q_reg_27 ( .CK(DNT_DW0_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW0[27]) );
    zdffqrb DNT_DW0_Q_reg_26 ( .CK(DNT_DW0_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW0[26]) );
    zdffqrb DNT_DW0_Q_reg_25 ( .CK(DNT_DW0_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW0[25]) );
    zdffqrb DNT_DW0_Q_reg_24 ( .CK(DNT_DW0_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW0[24]) );
    zdffqrb DNT_DW0_Q_reg_23 ( .CK(DNT_DW0_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW0[23]) );
    zdffqrb DNT_DW0_Q_reg_22 ( .CK(DNT_DW0_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW0[22]) );
    zdffqrb DNT_DW0_Q_reg_21 ( .CK(DNT_DW0_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW0[21]) );
    zdffqrb DNT_DW0_Q_reg_20 ( .CK(DNT_DW0_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW0[20]) );
    zdffqrb DNT_DW0_Q_reg_19 ( .CK(DNT_DW0_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW0[19]) );
    zdffqrb DNT_DW0_Q_reg_18 ( .CK(DNT_DW0_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW0[18]) );
    zdffqrb DNT_DW0_Q_reg_17 ( .CK(DNT_DW0_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW0[17]) );
    zdffqrb DNT_DW0_Q_reg_16 ( .CK(DNT_DW0_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW0[16]) );
    zdffqrb DNT_DW0_Q_reg_15 ( .CK(DNT_DW0_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW0[15]) );
    zdffqrb DNT_DW0_Q_reg_14 ( .CK(DNT_DW0_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW0[14]) );
    zdffqrb DNT_DW0_Q_reg_13 ( .CK(DNT_DW0_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW0[13]) );
    zdffqrb DNT_DW0_Q_reg_12 ( .CK(DNT_DW0_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW0[12]) );
    zdffqrb DNT_DW0_Q_reg_11 ( .CK(DNT_DW0_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW0[11]) );
    zdffqrb DNT_DW0_Q_reg_10 ( .CK(DNT_DW0_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW0[10]) );
    zdffqrb DNT_DW0_Q_reg_9 ( .CK(DNT_DW0_n126), .D(ADI[9]), .R(TRST_), .Q(DW0
        [9]) );
    zdffqrb DNT_DW0_Q_reg_8 ( .CK(DNT_DW0_n126), .D(ADI[8]), .R(TRST_), .Q(DW0
        [8]) );
    zdffqrb DNT_DW0_Q_reg_7 ( .CK(DNT_DW0_n126), .D(ADI[7]), .R(TRST_), .Q(DW0
        [7]) );
    zdffqrb DNT_DW0_Q_reg_6 ( .CK(DNT_DW0_n126), .D(ADI[6]), .R(TRST_), .Q(DW0
        [6]) );
    zdffqrb DNT_DW0_Q_reg_5 ( .CK(DNT_DW0_n126), .D(ADI[5]), .R(TRST_), .Q(DW0
        [5]) );
    zdffqrb DNT_DW0_Q_reg_4 ( .CK(DNT_DW0_n126), .D(ADI[4]), .R(TRST_), .Q(DW0
        [4]) );
    zdffqrb DNT_DW0_Q_reg_3 ( .CK(DNT_DW0_n126), .D(ADI[3]), .R(TRST_), .Q(DW0
        [3]) );
    zdffqrb DNT_DW0_Q_reg_2 ( .CK(DNT_DW0_n126), .D(ADI[2]), .R(TRST_), .Q(DW0
        [2]) );
    zdffqrb DNT_DW0_Q_reg_1 ( .CK(DNT_DW0_n126), .D(ADI[1]), .R(TRST_), .Q(DW0
        [1]) );
    zdffqrb DNT_DW0_Q_reg_0 ( .CK(DNT_DW0_n126), .D(ADI[0]), .R(TRST_), .Q(DW0
        [0]) );
    zbfb DNT_DW0_U80 ( .A(FLOPS_CLK_14), .Y(DNT_DW0_n126) );
    zbfb DNT_DW0_U81 ( .A(FLOPS_CLK_14), .Y(DNT_DW0_n127) );
endmodule


module PERIODIC_CACHE ( LDW, ADI, PCICLK, TRST_, CACHE_EN, DW0, DW1, DW2, DW3, 
    DW4, DW5, DW6, DW7, DW8, DW9, DW10, DW11, DW12, DW13, DW14, DW15, 
    CACHEPHASE, UP_DW3, UP_DW4, UP_DW5, UP_DW6, UP_DW7, UP_DW8, UP_DW9, 
    UP_LDW3, UP_LDW4, UP_LDW5, UP_LDW6, UP_LDW7, UP_LDW8, UP_LDW9, ATPG_ENI );
input  [15:0] LDW;
output [31:0] DW0;
output [31:0] DW14;
input  [31:0] UP_DW8;
input  [31:0] ADI;
output [31:0] DW7;
output [31:0] DW9;
input  [31:0] UP_DW6;
output [31:0] DW13;
output [31:0] DW1;
output [31:0] DW6;
output [31:0] DW12;
input  [31:0] UP_DW7;
input  [31:0] UP_DW9;
output [31:0] DW2;
output [31:0] DW3;
output [31:0] DW8;
output [31:0] DW15;
output [31:0] DW4;
input  [31:0] UP_DW5;
output [31:0] DW5;
output [31:0] DW10;
output [31:0] DW11;
input  [31:0] UP_DW4;
input  [31:0] UP_DW3;
input  PCICLK, TRST_, CACHE_EN, CACHEPHASE, UP_LDW3, UP_LDW4, UP_LDW5, UP_LDW6, 
    UP_LDW7, UP_LDW8, UP_LDW9, ATPG_ENI;
    wire AD8IN_0, AD5IN_3, FLOPS_CLK_13, FLOPS_CLK_7, AD6IN_9, AD3IN_25, 
        AD8IN_14, AD9IN_26, AD3IN_2, AD7IN_21, AD7IN_5, AD6IN_13, AD5IN_10, 
        AD3IN_19, AD4IN_22, AD8IN_28, AD8IN_9, n_23, AD6IN_0, AD4IN_17, 
        AD9IN_5, AD4IN_30, AD4IN_6, AD5IN_25, n_7, AD7IN_28, AD6IN_26, 
        AD7IN_14, AD5IN_19, n_18, AD3IN_10, AD8IN_21, AD9IN_13, AD3IN_30, 
        AD3IN_17, AD8IN_26, AD9IN_14, AD7IN_13, AD6IN_21, AD4IN_1, AD5IN_22, 
        AD4IN_10, AD9IN_2, n_9, n_24, AD6IN_7, FLOPS_CLK_9, AD9IN_28, AD6IN_28, 
        AD4IN_25, AD5IN_30, AD5IN_17, AD4IN_19, AD3IN_5, AD4IN_8, AD6IN_14, 
        AD7IN_2, AD7IN_26, AD5IN_4, FLOPS_CLK_14, AD8IN_7, AD9IN_21, AD3IN_22, 
        AD8IN_13, FLOPS_CLK_0, AD6IN_6, AD4IN_0, AD9IN_29, FLOPS_CLK_8, 
        AD5IN_23, AD4IN_11, AD9IN_3, n_19, n_25, AD7IN_12, AD6IN_20, AD3IN_31, 
        AD3IN_16, AD8IN_27, AD9IN_15, FLOPS_CLK_15, AD5IN_5, AD8IN_6, n_8, 
        n_10, AD3IN_23, AD8IN_12, AD9IN_20, FLOPS_CLK_1, AD3IN_4, AD4IN_18, 
        AD4IN_9, AD6IN_15, AD7IN_3, AD7IN_27, AD6IN_29, AD4IN_24, AD5IN_31, 
        AD5IN_16, AD3IN_18, AD8IN_29, AD5IN_11, AD4IN_23, AD3IN_3, AD7IN_20, 
        AD7IN_4, AD6IN_12, AD8IN_1, AD5IN_2, AD6IN_8, FLOPS_CLK_12, AD3IN_24, 
        FLOPS_CLK_6, AD8IN_15, AD9IN_27, n_6, AD3IN_11, AD9IN_12, AD8IN_20, 
        AD6IN_27, AD7IN_15, n_22, AD5IN_18, AD4IN_16, AD9IN_4, AD4IN_31, 
        AD4IN_7, AD5IN_24, AD7IN_29, AD8IN_8, AD6IN_1, AD8IN_30, AD9IN_25, 
        FLOPS_CLK_4, AD3IN_26, AD8IN_17, AD5IN_0, FLOPS_CLK_10, AD7IN_6, 
        AD8IN_3, AD6IN_10, AD7IN_22, AD3IN_1, AD4IN_21, AD5IN_13, n_20, 
        AD6IN_3, AD9IN_19, AD5IN_9, AD6IN_19, AD3IN_8, AD4IN_14, AD4IN_5, 
        AD5IN_26, AD9IN_6, AD4IN_28, AD7IN_17, AD6IN_25, AD7IN_30, AD3IN_13, 
        AD8IN_22, AD9IN_10, AD9IN_17, AD3IN_14, AD9IN_30, AD8IN_25, n_27, 
        AD6IN_22, AD7IN_10, AD7IN_8, AD4IN_13, AD9IN_1, AD4IN_2, AD5IN_21, 
        AD3IN_28, AD6IN_4, AD8IN_19, AD4IN_26, AD5IN_14, AD7IN_19, AD6IN_30, 
        AD7IN_25, AD6IN_17, AD7IN_1, AD5IN_28, AD3IN_21, AD3IN_6, AD9IN_8, 
        AD8IN_10, FLOPS_CLK_3, AD9IN_22, n_26, AD8IN_4, AD5IN_7, AD3IN_29, 
        AD6IN_5, AD8IN_18, AD7IN_9, AD4IN_12, AD4IN_3, AD9IN_0, AD5IN_20, 
        AD6IN_23, AD7IN_11, AD9IN_16, AD3IN_20, AD3IN_15, AD8IN_24, AD9IN_31, 
        AD8IN_11, FLOPS_CLK_2, AD9IN_23, AD8IN_5, AD5IN_6, AD6IN_31, AD7IN_24, 
        AD6IN_16, AD7IN_0, AD5IN_29, AD3IN_7, AD9IN_9, AD4IN_27, AD5IN_15, 
        AD7IN_18, AD9IN_18, AD4IN_20, AD5IN_12, AD7IN_7, AD6IN_11, AD7IN_23, 
        AD3IN_0, AD8IN_31, AD9IN_24, AD3IN_27, FLOPS_CLK_5, AD5IN_1, AD8IN_16, 
        FLOPS_CLK_11, AD8IN_2, AD3IN_12, AD8IN_23, n_5, AD9IN_11, n_21, 
        AD4IN_29, AD7IN_16, AD6IN_24, AD7IN_31, AD6IN_18, AD3IN_9, AD4IN_4, 
        AD5IN_27, AD4IN_15, AD9IN_7, AD6IN_2, AD5IN_8, n410, n411, n412, n413, 
        n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
        n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
        n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, 
        n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, 
        n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, 
        n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, 
        n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, 
        n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
        DNT_DW6_n126, DNT_DW6_n127, DNT_DW1_n126, DNT_DW1_n127, DNT_DW10_n126, 
        DNT_DW10_n127, DNT_DW8_n126, DNT_DW8_n127, DNT_DW0_n126, DNT_DW0_n127, 
        DNT_DW11_n126, DNT_DW11_n127, DNT_DW9_n126, DNT_DW9_n127, DNT_DW7_n126, 
        DNT_DW7_n127, DNT_DW5_n126, DNT_DW5_n127, DNT_DW14_n126, DNT_DW14_n127, 
        DNT_DW2_n126, DNT_DW2_n127, DNT_DW13_n126, DNT_DW13_n127, DNT_DW3_n126, 
        DNT_DW3_n127, DNT_DW12_n126, DNT_DW12_n127, DNT_DW4_n126, DNT_DW4_n127, 
        DNT_DW15_n126, DNT_DW15_n127;
    zan2b U61 ( .A(LDW[15]), .B(n442), .Y(n_5) );
    zao21b U62 ( .A(LDW[4]), .B(CACHE_EN), .C(UP_LDW4), .Y(n_26) );
    zan2b U63 ( .A(LDW[12]), .B(n442), .Y(n_8) );
    zao21b U64 ( .A(LDW[3]), .B(CACHE_EN), .C(UP_LDW3), .Y(n_27) );
    zan2b U65 ( .A(LDW[13]), .B(n442), .Y(n_7) );
    zan2b U66 ( .A(LDW[2]), .B(n442), .Y(n_18) );
    zan2b U67 ( .A(LDW[14]), .B(n442), .Y(n_6) );
    zao21b U68 ( .A(LDW[5]), .B(CACHE_EN), .C(UP_LDW5), .Y(n_25) );
    zao21b U69 ( .A(LDW[7]), .B(CACHE_EN), .C(UP_LDW7), .Y(n_23) );
    zao21b U70 ( .A(LDW[9]), .B(CACHE_EN), .C(UP_LDW9), .Y(n_21) );
    zan2b U71 ( .A(n442), .B(LDW[11]), .Y(n_9) );
    zan2b U72 ( .A(LDW[0]), .B(n442), .Y(n_20) );
    zao21b U73 ( .A(LDW[8]), .B(CACHE_EN), .C(UP_LDW8), .Y(n_22) );
    zan2b U74 ( .A(LDW[10]), .B(n442), .Y(n_10) );
    zan2b U75 ( .A(LDW[1]), .B(n442), .Y(n_19) );
    zbfb U76 ( .A(CACHE_EN), .Y(n442) );
    zao21b U77 ( .A(LDW[6]), .B(CACHE_EN), .C(UP_LDW6), .Y(n_24) );
    zao21b U78 ( .A(UP_DW4[1]), .B(n496), .C(n440), .Y(AD4IN_1) );
    zao21b U79 ( .A(UP_DW4[4]), .B(n498), .C(n437), .Y(AD4IN_4) );
    zao21b U80 ( .A(UP_DW4[6]), .B(n500), .C(n435), .Y(AD4IN_6) );
    zao21b U81 ( .A(UP_DW4[8]), .B(n481), .C(n433), .Y(AD4IN_8) );
    zao21b U82 ( .A(UP_DW4[10]), .B(n482), .C(n431), .Y(AD4IN_10) );
    zao21b U83 ( .A(UP_DW4[14]), .B(n481), .C(n427), .Y(AD4IN_14) );
    zao21b U84 ( .A(UP_DW4[16]), .B(n496), .C(n425), .Y(AD4IN_16) );
    zao21b U85 ( .A(UP_DW4[18]), .B(n491), .C(n423), .Y(AD4IN_18) );
    zao21b U86 ( .A(UP_DW4[20]), .B(n506), .C(n421), .Y(AD4IN_20) );
    zao21b U87 ( .A(UP_DW4[22]), .B(n496), .C(n419), .Y(AD4IN_22) );
    zao21b U88 ( .A(UP_DW4[26]), .B(n503), .C(n415), .Y(AD4IN_26) );
    zao21b U89 ( .A(UP_DW3[0]), .B(n506), .C(n441), .Y(AD3IN_0) );
    zao21b U90 ( .A(UP_DW3[3]), .B(n487), .C(n438), .Y(AD3IN_3) );
    zao21b U91 ( .A(UP_DW3[7]), .B(n493), .C(n434), .Y(AD3IN_7) );
    zao21b U92 ( .A(UP_DW3[8]), .B(n483), .C(n433), .Y(AD3IN_8) );
    zao21b U93 ( .A(UP_DW3[12]), .B(n495), .C(n429), .Y(AD3IN_12) );
    zao21b U94 ( .A(UP_DW3[17]), .B(n478), .C(n424), .Y(AD3IN_17) );
    zao21b U95 ( .A(UP_DW3[18]), .B(n490), .C(n423), .Y(AD3IN_18) );
    zao21b U96 ( .A(UP_DW3[19]), .B(n488), .C(n422), .Y(AD3IN_19) );
    zao21b U97 ( .A(UP_DW3[20]), .B(n478), .C(n421), .Y(AD3IN_20) );
    zao21b U98 ( .A(UP_DW3[23]), .B(n497), .C(n418), .Y(AD3IN_23) );
    zao21b U99 ( .A(UP_DW3[26]), .B(n498), .C(n415), .Y(AD3IN_26) );
    zao21b U100 ( .A(UP_DW3[27]), .B(n503), .C(n414), .Y(AD3IN_27) );
    zao21b U101 ( .A(UP_DW5[0]), .B(n504), .C(n441), .Y(AD5IN_0) );
    zao21b U102 ( .A(UP_DW5[1]), .B(n497), .C(n440), .Y(AD5IN_1) );
    zao21b U103 ( .A(UP_DW5[3]), .B(n482), .C(n438), .Y(AD5IN_3) );
    zao21b U104 ( .A(UP_DW5[4]), .B(n477), .C(n437), .Y(AD5IN_4) );
    zao21b U105 ( .A(UP_DW5[5]), .B(n443), .C(n436), .Y(AD5IN_5) );
    zao21b U106 ( .A(UP_DW5[6]), .B(n480), .C(n435), .Y(AD5IN_6) );
    zao21b U107 ( .A(UP_DW5[10]), .B(n489), .C(n431), .Y(AD5IN_10) );
    zao21b U108 ( .A(UP_DW5[11]), .B(n485), .C(n430), .Y(AD5IN_11) );
    zao21b U109 ( .A(UP_DW5[13]), .B(n496), .C(n428), .Y(AD5IN_13) );
    zao21b U110 ( .A(UP_DW5[14]), .B(n500), .C(n427), .Y(AD5IN_14) );
    zao21b U111 ( .A(UP_DW5[15]), .B(n481), .C(n426), .Y(AD5IN_15) );
    zao21b U112 ( .A(UP_DW5[16]), .B(n477), .C(n425), .Y(AD5IN_16) );
    zao21b U113 ( .A(UP_DW5[21]), .B(n497), .C(n420), .Y(AD5IN_21) );
    zao21b U114 ( .A(UP_DW5[22]), .B(n489), .C(n419), .Y(AD5IN_22) );
    zao21b U115 ( .A(UP_DW5[23]), .B(n503), .C(n418), .Y(AD5IN_23) );
    zao21b U116 ( .A(UP_DW5[24]), .B(n443), .C(n417), .Y(AD5IN_24) );
    zao21b U117 ( .A(UP_DW5[25]), .B(n477), .C(n416), .Y(AD5IN_25) );
    zao21b U118 ( .A(UP_DW5[26]), .B(n486), .C(n415), .Y(AD5IN_26) );
    zao21b U119 ( .A(UP_DW5[28]), .B(n497), .C(n413), .Y(AD5IN_28) );
    zao21b U120 ( .A(UP_DW5[29]), .B(n478), .C(n412), .Y(AD5IN_29) );
    zao21b U121 ( .A(UP_DW5[30]), .B(n501), .C(n411), .Y(AD5IN_30) );
    zao21b U122 ( .A(UP_DW5[31]), .B(n496), .C(n410), .Y(AD5IN_31) );
    zao21b U123 ( .A(UP_DW7[7]), .B(n489), .C(n434), .Y(AD7IN_7) );
    zao21b U124 ( .A(UP_DW7[9]), .B(n486), .C(n432), .Y(AD7IN_9) );
    zao21b U125 ( .A(UP_DW7[11]), .B(n484), .C(n430), .Y(AD7IN_11) );
    zao21b U126 ( .A(UP_DW7[12]), .B(n486), .C(n429), .Y(AD7IN_12) );
    zao21b U127 ( .A(UP_DW7[13]), .B(n498), .C(n428), .Y(AD7IN_13) );
    zao21b U128 ( .A(UP_DW7[16]), .B(n489), .C(n425), .Y(AD7IN_16) );
    zao21b U129 ( .A(UP_DW7[18]), .B(n495), .C(n423), .Y(AD7IN_18) );
    zao21b U130 ( .A(UP_DW7[20]), .B(n485), .C(n421), .Y(AD7IN_20) );
    zao21b U131 ( .A(UP_DW7[21]), .B(n491), .C(n420), .Y(AD7IN_21) );
    zao21b U132 ( .A(UP_DW7[22]), .B(n504), .C(n419), .Y(AD7IN_22) );
    zao21b U133 ( .A(UP_DW7[23]), .B(n481), .C(n418), .Y(AD7IN_23) );
    zao21b U134 ( .A(UP_DW7[24]), .B(n504), .C(n417), .Y(AD7IN_24) );
    zao21b U135 ( .A(UP_DW7[26]), .B(n500), .C(n415), .Y(AD7IN_26) );
    zao21b U136 ( .A(UP_DW7[27]), .B(n491), .C(n414), .Y(AD7IN_27) );
    zao21b U137 ( .A(UP_DW7[30]), .B(n477), .C(n411), .Y(AD7IN_30) );
    zao21b U138 ( .A(UP_DW7[31]), .B(n480), .C(n410), .Y(AD7IN_31) );
    zao21b U139 ( .A(UP_DW9[4]), .B(n495), .C(n437), .Y(AD9IN_4) );
    zao21b U140 ( .A(UP_DW9[5]), .B(n487), .C(n436), .Y(AD9IN_5) );
    zao21b U141 ( .A(UP_DW9[6]), .B(n492), .C(n435), .Y(AD9IN_6) );
    zao21b U142 ( .A(n504), .B(UP_DW9[9]), .C(n432), .Y(AD9IN_9) );
    zao21b U143 ( .A(UP_DW9[11]), .B(n482), .C(n430), .Y(AD9IN_11) );
    zao21b U144 ( .A(UP_DW9[12]), .B(n488), .C(n429), .Y(AD9IN_12) );
    zao21b U145 ( .A(UP_DW9[19]), .B(n492), .C(n422), .Y(AD9IN_19) );
    zao21b U146 ( .A(UP_DW9[20]), .B(n503), .C(n421), .Y(AD9IN_20) );
    zao21b U147 ( .A(UP_DW9[22]), .B(n484), .C(n419), .Y(AD9IN_22) );
    zao21b U148 ( .A(UP_DW9[23]), .B(n488), .C(n418), .Y(AD9IN_23) );
    zao21b U149 ( .A(UP_DW9[24]), .B(n483), .C(n417), .Y(AD9IN_24) );
    zao21b U150 ( .A(UP_DW9[26]), .B(n505), .C(n415), .Y(AD9IN_26) );
    zao21b U151 ( .A(UP_DW9[27]), .B(n487), .C(n414), .Y(AD9IN_27) );
    zao21b U152 ( .A(UP_DW9[29]), .B(n498), .C(n412), .Y(AD9IN_29) );
    zao21b U153 ( .A(UP_DW9[31]), .B(n443), .C(n410), .Y(AD9IN_31) );
    zao21b U154 ( .A(UP_DW8[1]), .B(n505), .C(n440), .Y(AD8IN_1) );
    zao21b U155 ( .A(UP_DW8[2]), .B(n498), .C(n439), .Y(AD8IN_2) );
    zao21b U156 ( .A(UP_DW8[5]), .B(n505), .C(n436), .Y(AD8IN_5) );
    zao21b U157 ( .A(UP_DW8[6]), .B(n486), .C(n435), .Y(AD8IN_6) );
    zao21b U158 ( .A(UP_DW8[7]), .B(n487), .C(n434), .Y(AD8IN_7) );
    zao21b U159 ( .A(UP_DW8[8]), .B(n506), .C(n433), .Y(AD8IN_8) );
    zao21b U160 ( .A(UP_DW8[11]), .B(n504), .C(n430), .Y(AD8IN_11) );
    zao21b U161 ( .A(UP_DW8[19]), .B(n443), .C(n422), .Y(AD8IN_19) );
    zao21b U162 ( .A(UP_DW8[21]), .B(n483), .C(n420), .Y(AD8IN_21) );
    zao21b U163 ( .A(UP_DW8[22]), .B(n491), .C(n419), .Y(AD8IN_22) );
    zao21b U164 ( .A(UP_DW8[23]), .B(n506), .C(n418), .Y(AD8IN_23) );
    zao21b U165 ( .A(UP_DW8[26]), .B(n483), .C(n415), .Y(AD8IN_26) );
    zao21b U166 ( .A(UP_DW6[1]), .B(n487), .C(n440), .Y(AD6IN_1) );
    zao21b U167 ( .A(UP_DW6[3]), .B(n488), .C(n438), .Y(AD6IN_3) );
    zao21b U168 ( .A(UP_DW6[4]), .B(n478), .C(n437), .Y(AD6IN_4) );
    zao21b U169 ( .A(UP_DW6[9]), .B(n482), .C(n432), .Y(AD6IN_9) );
    zao21b U170 ( .A(UP_DW6[10]), .B(n480), .C(n431), .Y(AD6IN_10) );
    zao21b U171 ( .A(UP_DW6[11]), .B(n500), .C(n430), .Y(AD6IN_11) );
    zao21b U172 ( .A(UP_DW6[15]), .B(n477), .C(n426), .Y(AD6IN_15) );
    zao21b U173 ( .A(UP_DW6[16]), .B(n480), .C(n425), .Y(AD6IN_16) );
    zao21b U174 ( .A(UP_DW6[18]), .B(n488), .C(n423), .Y(AD6IN_18) );
    zao21b U175 ( .A(UP_DW6[19]), .B(n505), .C(n422), .Y(AD6IN_19) );
    zao21b U176 ( .A(UP_DW6[22]), .B(n480), .C(n419), .Y(AD6IN_22) );
    zao21b U177 ( .A(UP_DW6[25]), .B(n486), .C(n416), .Y(AD6IN_25) );
    zao21b U178 ( .A(UP_DW6[26]), .B(n443), .C(n415), .Y(AD6IN_26) );
    zao21b U179 ( .A(UP_DW6[27]), .B(n483), .C(n414), .Y(AD6IN_27) );
    zao21b U180 ( .A(UP_DW6[28]), .B(n478), .C(n413), .Y(AD6IN_28) );
    zao21b U181 ( .A(UP_DW6[29]), .B(n501), .C(n412), .Y(AD6IN_29) );
    zao21b U182 ( .A(UP_DW6[30]), .B(n495), .C(n411), .Y(AD6IN_30) );
    zao21b U183 ( .A(UP_DW6[31]), .B(n505), .C(n410), .Y(AD6IN_31) );
    zan2b U184 ( .A(ADI[31]), .B(n479), .Y(n410) );
    zan2b U185 ( .A(ADI[30]), .B(n507), .Y(n411) );
    zan2b U186 ( .A(ADI[29]), .B(n508), .Y(n412) );
    zan2b U187 ( .A(ADI[28]), .B(n479), .Y(n413) );
    zan2b U188 ( .A(ADI[27]), .B(n507), .Y(n414) );
    zan2b U189 ( .A(ADI[26]), .B(n444), .Y(n415) );
    zan2b U190 ( .A(ADI[25]), .B(n508), .Y(n416) );
    zan2b U191 ( .A(ADI[24]), .B(n479), .Y(n417) );
    zan2b U192 ( .A(ADI[23]), .B(n444), .Y(n418) );
    zan2b U193 ( .A(ADI[22]), .B(n507), .Y(n419) );
    zan2b U194 ( .A(ADI[21]), .B(n479), .Y(n420) );
    zan2b U195 ( .A(ADI[20]), .B(n508), .Y(n421) );
    zan2b U196 ( .A(ADI[19]), .B(n444), .Y(n422) );
    zan2b U197 ( .A(ADI[18]), .B(n444), .Y(n423) );
    zan2b U198 ( .A(ADI[17]), .B(n444), .Y(n424) );
    zan2b U199 ( .A(ADI[16]), .B(n508), .Y(n425) );
    zan2b U200 ( .A(ADI[15]), .B(n507), .Y(n426) );
    zan2b U201 ( .A(ADI[14]), .B(n479), .Y(n427) );
    zan2b U202 ( .A(ADI[13]), .B(n508), .Y(n428) );
    zan2b U203 ( .A(ADI[12]), .B(n479), .Y(n429) );
    zan2b U204 ( .A(ADI[11]), .B(n508), .Y(n430) );
    zan2b U205 ( .A(ADI[10]), .B(n444), .Y(n431) );
    zan2b U206 ( .A(ADI[9]), .B(n507), .Y(n432) );
    zan2b U207 ( .A(ADI[8]), .B(n508), .Y(n433) );
    zan2b U208 ( .A(ADI[7]), .B(n444), .Y(n434) );
    zan2b U209 ( .A(ADI[6]), .B(n444), .Y(n435) );
    zan2b U210 ( .A(ADI[5]), .B(n508), .Y(n436) );
    zan2b U211 ( .A(ADI[4]), .B(n507), .Y(n437) );
    zan2b U212 ( .A(ADI[3]), .B(n444), .Y(n438) );
    zan2b U213 ( .A(ADI[2]), .B(n507), .Y(n439) );
    zan2b U214 ( .A(ADI[1]), .B(n508), .Y(n440) );
    zan2b U215 ( .A(ADI[0]), .B(n507), .Y(n441) );
    ziv11b U216 ( .A(n499), .Y(n443), .Z(n444) );
    zbfb U217 ( .A(ADI[31]), .Y(n445) );
    zbfb U218 ( .A(ADI[16]), .Y(n446) );
    zbfb U219 ( .A(ADI[7]), .Y(n447) );
    zbfb U220 ( .A(ADI[11]), .Y(n448) );
    zbfb U221 ( .A(ADI[23]), .Y(n449) );
    zbfb U222 ( .A(ADI[0]), .Y(n450) );
    zbfb U223 ( .A(ADI[5]), .Y(n451) );
    zbfb U224 ( .A(ADI[18]), .Y(n452) );
    zbfb U225 ( .A(ADI[28]), .Y(n453) );
    zbfb U226 ( .A(ADI[9]), .Y(n454) );
    zbfb U227 ( .A(ADI[14]), .Y(n455) );
    zbfb U228 ( .A(ADI[24]), .Y(n456) );
    zbfb U229 ( .A(ADI[21]), .Y(n457) );
    zbfb U230 ( .A(ADI[1]), .Y(n458) );
    zbfb U231 ( .A(ADI[26]), .Y(n459) );
    zbfb U232 ( .A(ADI[10]), .Y(n460) );
    zbfb U233 ( .A(ADI[13]), .Y(n461) );
    zbfb U234 ( .A(ADI[8]), .Y(n462) );
    zbfb U235 ( .A(ADI[2]), .Y(n463) );
    zbfb U236 ( .A(ADI[25]), .Y(n464) );
    zbfb U237 ( .A(ADI[27]), .Y(n465) );
    zbfb U238 ( .A(ADI[19]), .Y(n466) );
    zbfb U239 ( .A(ADI[3]), .Y(n467) );
    zbfb U240 ( .A(ADI[22]), .Y(n468) );
    zbfb U241 ( .A(ADI[12]), .Y(n469) );
    zbfb U242 ( .A(ADI[30]), .Y(n470) );
    zbfb U243 ( .A(ADI[15]), .Y(n471) );
    zbfb U244 ( .A(ADI[17]), .Y(n472) );
    zbfb U245 ( .A(ADI[4]), .Y(n473) );
    zbfb U246 ( .A(ADI[6]), .Y(n474) );
    zbfb U247 ( .A(ADI[29]), .Y(n475) );
    zbfb U248 ( .A(ADI[20]), .Y(n476) );
    zivb U249 ( .A(n494), .Y(n477) );
    zao21b U250 ( .A(UP_DW7[6]), .B(n489), .C(n435), .Y(AD7IN_6) );
    zao21b U251 ( .A(UP_DW7[29]), .B(n482), .C(n412), .Y(AD7IN_29) );
    zao21b U252 ( .A(UP_DW9[18]), .B(n497), .C(n423), .Y(AD9IN_18) );
    zao21b U253 ( .A(UP_DW8[24]), .B(n495), .C(n417), .Y(AD8IN_24) );
    zao21b U254 ( .A(UP_DW8[15]), .B(n498), .C(n426), .Y(AD8IN_15) );
    zao21b U255 ( .A(UP_DW5[17]), .B(n488), .C(n424), .Y(AD5IN_17) );
    zivb U256 ( .A(n502), .Y(n478) );
    zao21b U257 ( .A(UP_DW6[7]), .B(n504), .C(n434), .Y(AD6IN_7) );
    zao21b U258 ( .A(UP_DW9[15]), .B(n503), .C(n426), .Y(AD9IN_15) );
    zao21b U259 ( .A(UP_DW7[15]), .B(n506), .C(n426), .Y(AD7IN_15) );
    zao21b U260 ( .A(UP_DW3[30]), .B(n481), .C(n411), .Y(AD3IN_30) );
    zao21b U261 ( .A(UP_DW8[18]), .B(n487), .C(n423), .Y(AD8IN_18) );
    zao21b U262 ( .A(UP_DW8[29]), .B(n505), .C(n412), .Y(AD8IN_29) );
    zivb U263 ( .A(n443), .Y(n479) );
    zivb U264 ( .A(n502), .Y(n480) );
    zivb U265 ( .A(n502), .Y(n481) );
    zao21b U266 ( .A(UP_DW7[4]), .B(n503), .C(n437), .Y(AD7IN_4) );
    zao21b U267 ( .A(UP_DW8[30]), .B(n478), .C(n411), .Y(AD8IN_30) );
    zao21b U268 ( .A(UP_DW3[24]), .B(n504), .C(n417), .Y(AD3IN_24) );
    zao21b U269 ( .A(UP_DW3[21]), .B(n486), .C(n420), .Y(AD3IN_21) );
    zao21b U270 ( .A(UP_DW3[14]), .B(n503), .C(n427), .Y(AD3IN_14) );
    zao21b U271 ( .A(UP_DW7[28]), .B(n478), .C(n413), .Y(AD7IN_28) );
    zao21b U272 ( .A(UP_DW3[6]), .B(n506), .C(n435), .Y(AD3IN_6) );
    zao21b U273 ( .A(UP_DW3[9]), .B(n478), .C(n432), .Y(AD3IN_9) );
    zao21b U274 ( .A(UP_DW4[2]), .B(n506), .C(n439), .Y(AD4IN_2) );
    zivb U275 ( .A(n494), .Y(n483) );
    zivb U276 ( .A(n494), .Y(n482) );
    zao21b U277 ( .A(UP_DW7[1]), .B(n497), .C(n440), .Y(AD7IN_1) );
    zao21b U278 ( .A(UP_DW8[20]), .B(n495), .C(n421), .Y(AD8IN_20) );
    zao21b U279 ( .A(UP_DW3[16]), .B(n496), .C(n425), .Y(AD3IN_16) );
    zao21b U280 ( .A(UP_DW4[25]), .B(n496), .C(n416), .Y(AD4IN_25) );
    zao21b U281 ( .A(UP_DW8[12]), .B(n489), .C(n429), .Y(AD8IN_12) );
    zao21b U282 ( .A(UP_DW9[30]), .B(n477), .C(n411), .Y(AD9IN_30) );
    zao21b U283 ( .A(UP_DW6[6]), .B(n477), .C(n435), .Y(AD6IN_6) );
    zao21b U284 ( .A(UP_DW6[24]), .B(n477), .C(n417), .Y(AD6IN_24) );
    zao21b U285 ( .A(UP_DW4[13]), .B(n488), .C(n428), .Y(AD4IN_13) );
    zivb U286 ( .A(n499), .Y(n485) );
    zivb U287 ( .A(n499), .Y(n484) );
    zivb U288 ( .A(n502), .Y(n487) );
    zivb U289 ( .A(n502), .Y(n486) );
    zao21b U290 ( .A(UP_DW9[21]), .B(n503), .C(n420), .Y(AD9IN_21) );
    zao21b U291 ( .A(UP_DW5[12]), .B(n506), .C(n429), .Y(AD5IN_12) );
    zao21b U292 ( .A(UP_DW9[14]), .B(n486), .C(n427), .Y(AD9IN_14) );
    zao21b U293 ( .A(UP_DW9[2]), .B(n504), .C(n439), .Y(AD9IN_2) );
    zao21b U294 ( .A(UP_DW8[3]), .B(n481), .C(n438), .Y(AD8IN_3) );
    zao21b U295 ( .A(UP_DW7[10]), .B(n504), .C(n431), .Y(AD7IN_10) );
    zao21b U296 ( .A(UP_DW6[13]), .B(n487), .C(n428), .Y(AD6IN_13) );
    zao21b U297 ( .A(UP_DW7[0]), .B(n487), .C(n441), .Y(AD7IN_0) );
    zao21b U298 ( .A(UP_DW9[17]), .B(n480), .C(n424), .Y(AD9IN_17) );
    zao21b U299 ( .A(UP_DW5[7]), .B(n480), .C(n434), .Y(AD5IN_7) );
    zao21b U300 ( .A(UP_DW7[3]), .B(n481), .C(n438), .Y(AD7IN_3) );
    zao21b U301 ( .A(UP_DW4[17]), .B(n480), .C(n424), .Y(AD4IN_17) );
    zao21b U302 ( .A(UP_DW4[5]), .B(n487), .C(n436), .Y(AD4IN_5) );
    zao21b U303 ( .A(UP_DW8[17]), .B(n505), .C(n424), .Y(AD8IN_17) );
    zao21b U304 ( .A(UP_DW5[9]), .B(n505), .C(n432), .Y(AD5IN_9) );
    zao21b U305 ( .A(UP_DW4[23]), .B(n505), .C(n418), .Y(AD4IN_23) );
    zao21b U306 ( .A(UP_DW4[29]), .B(n481), .C(n412), .Y(AD4IN_29) );
    zao21b U307 ( .A(UP_DW8[9]), .B(n486), .C(n432), .Y(AD8IN_9) );
    zao21b U308 ( .A(UP_DW4[11]), .B(n486), .C(n430), .Y(AD4IN_11) );
    zivb U309 ( .A(n494), .Y(n488) );
    zivb U310 ( .A(n494), .Y(n489) );
    zao21b U311 ( .A(UP_DW4[28]), .B(n488), .C(n413), .Y(AD4IN_28) );
    zao21b U312 ( .A(UP_DW7[19]), .B(n488), .C(n422), .Y(AD7IN_19) );
    zao21b U313 ( .A(UP_DW5[19]), .B(n498), .C(n422), .Y(AD5IN_19) );
    zao21b U314 ( .A(UP_DW8[0]), .B(n489), .C(n441), .Y(AD8IN_0) );
    zao21b U315 ( .A(UP_DW3[29]), .B(n498), .C(n412), .Y(AD3IN_29) );
    zao21b U316 ( .A(UP_DW9[8]), .B(n495), .C(n433), .Y(AD9IN_8) );
    zao21b U317 ( .A(UP_DW5[18]), .B(n477), .C(n423), .Y(AD5IN_18) );
    zao21b U318 ( .A(UP_DW9[10]), .B(n483), .C(n431), .Y(AD9IN_10) );
    zao21b U319 ( .A(UP_DW6[0]), .B(n483), .C(n441), .Y(AD6IN_0) );
    zao21b U320 ( .A(UP_DW8[14]), .B(n497), .C(n427), .Y(AD8IN_14) );
    zao21b U321 ( .A(UP_DW4[19]), .B(n495), .C(n422), .Y(AD4IN_19) );
    zao21b U322 ( .A(UP_DW8[27]), .B(n482), .C(n414), .Y(AD8IN_27) );
    zao21b U323 ( .A(UP_DW3[2]), .B(n498), .C(n439), .Y(AD3IN_2) );
    zao21b U324 ( .A(UP_DW9[3]), .B(n482), .C(n438), .Y(AD9IN_3) );
    zao21b U325 ( .A(UP_DW6[12]), .B(n489), .C(n429), .Y(AD6IN_12) );
    zao21b U326 ( .A(UP_DW6[21]), .B(n483), .C(n420), .Y(AD6IN_21) );
    zao21b U327 ( .A(UP_DW3[5]), .B(n496), .C(n436), .Y(AD3IN_5) );
    zao21b U328 ( .A(UP_DW5[20]), .B(n482), .C(n421), .Y(AD5IN_20) );
    zao21b U329 ( .A(UP_DW4[7]), .B(n497), .C(n434), .Y(AD4IN_7) );
    zivb U330 ( .A(n499), .Y(n491) );
    zivb U331 ( .A(n499), .Y(n490) );
    zao21b U332 ( .A(UP_DW9[7]), .B(n501), .C(n434), .Y(AD9IN_7) );
    zao21b U333 ( .A(UP_DW5[8]), .B(n501), .C(n433), .Y(AD5IN_8) );
    zao21b U334 ( .A(UP_DW4[12]), .B(n490), .C(n429), .Y(AD4IN_12) );
    zao21b U335 ( .A(UP_DW8[25]), .B(n501), .C(n416), .Y(AD8IN_25) );
    zao21b U336 ( .A(UP_DW9[25]), .B(n501), .C(n416), .Y(AD9IN_25) );
    zao21b U337 ( .A(UP_DW4[31]), .B(n484), .C(n410), .Y(AD4IN_31) );
    zao21b U338 ( .A(UP_DW6[23]), .B(n490), .C(n418), .Y(AD6IN_23) );
    zao21b U339 ( .A(UP_DW3[25]), .B(n490), .C(n416), .Y(AD3IN_25) );
    zao21b U340 ( .A(UP_DW6[14]), .B(n501), .C(n427), .Y(AD6IN_14) );
    zao21b U341 ( .A(UP_DW4[9]), .B(n492), .C(n432), .Y(AD4IN_9) );
    zao21b U342 ( .A(UP_DW7[25]), .B(n490), .C(n416), .Y(AD7IN_25) );
    zao21b U343 ( .A(UP_DW5[2]), .B(n490), .C(n439), .Y(AD5IN_2) );
    zao21b U344 ( .A(UP_DW3[28]), .B(n493), .C(n413), .Y(AD3IN_28) );
    zao21b U345 ( .A(UP_DW3[10]), .B(n493), .C(n431), .Y(AD3IN_10) );
    zao21b U346 ( .A(UP_DW8[13]), .B(n484), .C(n428), .Y(AD8IN_13) );
    zao21b U347 ( .A(UP_DW4[27]), .B(n484), .C(n414), .Y(AD4IN_27) );
    zao21b U348 ( .A(UP_DW7[14]), .B(n493), .C(n427), .Y(AD7IN_14) );
    zao21b U349 ( .A(UP_DW7[2]), .B(n492), .C(n439), .Y(AD7IN_2) );
    zao21b U350 ( .A(UP_DW6[2]), .B(n492), .C(n439), .Y(AD6IN_2) );
    zao21b U351 ( .A(UP_DW8[31]), .B(n484), .C(n410), .Y(AD8IN_31) );
    zao21b U352 ( .A(UP_DW9[1]), .B(n485), .C(n440), .Y(AD9IN_1) );
    zao21b U353 ( .A(UP_DW3[4]), .B(n490), .C(n437), .Y(AD3IN_4) );
    zao21b U354 ( .A(UP_DW4[0]), .B(n490), .C(n441), .Y(AD4IN_0) );
    zao21b U355 ( .A(UP_DW7[5]), .B(n493), .C(n436), .Y(AD7IN_5) );
    zivb U356 ( .A(n499), .Y(n500) );
    zivb U357 ( .A(n499), .Y(n492) );
    zivb U358 ( .A(n499), .Y(n493) );
    zao21b U359 ( .A(UP_DW9[28]), .B(n493), .C(n413), .Y(AD9IN_28) );
    zao21b U360 ( .A(UP_DW8[28]), .B(n493), .C(n413), .Y(AD8IN_28) );
    zao21b U361 ( .A(UP_DW6[5]), .B(n443), .C(n436), .Y(AD6IN_5) );
    zao21b U362 ( .A(UP_DW8[16]), .B(n485), .C(n425), .Y(AD8IN_16) );
    zao21b U363 ( .A(UP_DW7[17]), .B(n500), .C(n424), .Y(AD7IN_17) );
    zao21b U364 ( .A(UP_DW5[27]), .B(n491), .C(n414), .Y(AD5IN_27) );
    zao21b U365 ( .A(UP_DW4[3]), .B(n484), .C(n438), .Y(AD4IN_3) );
    zao21b U366 ( .A(UP_DW3[22]), .B(n500), .C(n419), .Y(AD3IN_22) );
    zao21b U367 ( .A(UP_DW6[17]), .B(n501), .C(n424), .Y(AD6IN_17) );
    zao21b U368 ( .A(UP_DW3[15]), .B(n492), .C(n426), .Y(AD3IN_15) );
    zao21b U369 ( .A(UP_DW3[13]), .B(n501), .C(n428), .Y(AD3IN_13) );
    zao21b U370 ( .A(UP_DW9[0]), .B(n492), .C(n441), .Y(AD9IN_0) );
    zao21b U371 ( .A(UP_DW8[4]), .B(n485), .C(n437), .Y(AD8IN_4) );
    zao21b U372 ( .A(UP_DW4[24]), .B(n493), .C(n417), .Y(AD4IN_24) );
    zao21b U373 ( .A(UP_DW3[11]), .B(n485), .C(n430), .Y(AD3IN_11) );
    zao21b U374 ( .A(UP_DW4[15]), .B(n484), .C(n426), .Y(AD4IN_15) );
    zao21b U375 ( .A(UP_DW6[20]), .B(n443), .C(n421), .Y(AD6IN_20) );
    zao21b U376 ( .A(UP_DW3[31]), .B(n493), .C(n410), .Y(AD3IN_31) );
    zao21b U377 ( .A(UP_DW4[30]), .B(n443), .C(n411), .Y(AD4IN_30) );
    zao21b U378 ( .A(UP_DW8[10]), .B(n484), .C(n431), .Y(AD8IN_10) );
    zao21b U379 ( .A(UP_DW3[1]), .B(n492), .C(n440), .Y(AD3IN_1) );
    zao21b U380 ( .A(UP_DW9[13]), .B(n485), .C(n428), .Y(AD9IN_13) );
    zao21b U381 ( .A(UP_DW7[8]), .B(n485), .C(n433), .Y(AD7IN_8) );
    zao21b U382 ( .A(UP_DW9[16]), .B(n485), .C(n425), .Y(AD9IN_16) );
    zao21b U383 ( .A(UP_DW4[21]), .B(n490), .C(n420), .Y(AD4IN_21) );
    zao21b U384 ( .A(UP_DW6[8]), .B(n492), .C(n433), .Y(AD6IN_8) );
    zivb U385 ( .A(n499), .Y(n501) );
    zivb U386 ( .A(CACHEPHASE), .Y(n494) );
    zivb U387 ( .A(n494), .Y(n495) );
    zivb U388 ( .A(n494), .Y(n498) );
    zivb U389 ( .A(n494), .Y(n496) );
    zivb U390 ( .A(n494), .Y(n497) );
    zivb U391 ( .A(CACHEPHASE), .Y(n499) );
    zivb U392 ( .A(n491), .Y(n508) );
    zivb U393 ( .A(n500), .Y(n507) );
    zivb U394 ( .A(CACHEPHASE), .Y(n502) );
    zivb U395 ( .A(n502), .Y(n503) );
    zivb U396 ( .A(n502), .Y(n506) );
    zivb U397 ( .A(n502), .Y(n504) );
    zivb U398 ( .A(n502), .Y(n505) );
    zmux21hd U399 ( .A(n_5), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_15) );
    zmux21hd U400 ( .A(n_6), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_14) );
    zmux21hd U401 ( .A(n_7), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_13) );
    zmux21hd U402 ( .A(n_8), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_12) );
    zmux21hd U403 ( .A(n_9), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_11) );
    zmux21hd U404 ( .A(n_10), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_10) );
    zmux21hd U405 ( .A(n_21), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_9) );
    zmux21hd U406 ( .A(n_22), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_8) );
    zmux21hd U407 ( .A(n_23), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_7) );
    zmux21hd U408 ( .A(n_24), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_6) );
    zmux21hd U409 ( .A(n_25), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_5) );
    zmux21hd U410 ( .A(n_26), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_4) );
    zmux21hd U411 ( .A(n_27), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_3) );
    zmux21hd U412 ( .A(n_18), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_2) );
    zmux21hd U413 ( .A(n_19), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_1) );
    zmux21hd U414 ( .A(n_20), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_0) );
    zdffqrb DNT_DW6_Q_reg_31 ( .CK(DNT_DW6_n127), .D(AD6IN_31), .R(TRST_), .Q(
        DW6[31]) );
    zdffqrb DNT_DW6_Q_reg_30 ( .CK(DNT_DW6_n127), .D(AD6IN_30), .R(TRST_), .Q(
        DW6[30]) );
    zdffqrb DNT_DW6_Q_reg_29 ( .CK(DNT_DW6_n127), .D(AD6IN_29), .R(TRST_), .Q(
        DW6[29]) );
    zdffqrb DNT_DW6_Q_reg_28 ( .CK(DNT_DW6_n127), .D(AD6IN_28), .R(TRST_), .Q(
        DW6[28]) );
    zdffqrb DNT_DW6_Q_reg_27 ( .CK(DNT_DW6_n127), .D(AD6IN_27), .R(TRST_), .Q(
        DW6[27]) );
    zdffqrb DNT_DW6_Q_reg_26 ( .CK(DNT_DW6_n127), .D(AD6IN_26), .R(TRST_), .Q(
        DW6[26]) );
    zdffqrb DNT_DW6_Q_reg_25 ( .CK(DNT_DW6_n127), .D(AD6IN_25), .R(TRST_), .Q(
        DW6[25]) );
    zdffqrb DNT_DW6_Q_reg_24 ( .CK(DNT_DW6_n127), .D(AD6IN_24), .R(TRST_), .Q(
        DW6[24]) );
    zdffqrb DNT_DW6_Q_reg_23 ( .CK(DNT_DW6_n127), .D(AD6IN_23), .R(TRST_), .Q(
        DW6[23]) );
    zdffqrb DNT_DW6_Q_reg_22 ( .CK(DNT_DW6_n127), .D(AD6IN_22), .R(TRST_), .Q(
        DW6[22]) );
    zdffqrb DNT_DW6_Q_reg_21 ( .CK(DNT_DW6_n127), .D(AD6IN_21), .R(TRST_), .Q(
        DW6[21]) );
    zdffqrb DNT_DW6_Q_reg_20 ( .CK(DNT_DW6_n127), .D(AD6IN_20), .R(TRST_), .Q(
        DW6[20]) );
    zdffqrb DNT_DW6_Q_reg_19 ( .CK(DNT_DW6_n127), .D(AD6IN_19), .R(TRST_), .Q(
        DW6[19]) );
    zdffqrb DNT_DW6_Q_reg_18 ( .CK(DNT_DW6_n127), .D(AD6IN_18), .R(TRST_), .Q(
        DW6[18]) );
    zdffqrb DNT_DW6_Q_reg_17 ( .CK(DNT_DW6_n127), .D(AD6IN_17), .R(TRST_), .Q(
        DW6[17]) );
    zdffqrb DNT_DW6_Q_reg_16 ( .CK(DNT_DW6_n127), .D(AD6IN_16), .R(TRST_), .Q(
        DW6[16]) );
    zdffqrb DNT_DW6_Q_reg_15 ( .CK(DNT_DW6_n126), .D(AD6IN_15), .R(TRST_), .Q(
        DW6[15]) );
    zdffqrb DNT_DW6_Q_reg_14 ( .CK(DNT_DW6_n126), .D(AD6IN_14), .R(TRST_), .Q(
        DW6[14]) );
    zdffqrb DNT_DW6_Q_reg_13 ( .CK(DNT_DW6_n126), .D(AD6IN_13), .R(TRST_), .Q(
        DW6[13]) );
    zdffqrb DNT_DW6_Q_reg_12 ( .CK(DNT_DW6_n126), .D(AD6IN_12), .R(TRST_), .Q(
        DW6[12]) );
    zdffqrb DNT_DW6_Q_reg_11 ( .CK(DNT_DW6_n126), .D(AD6IN_11), .R(TRST_), .Q(
        DW6[11]) );
    zdffqrb DNT_DW6_Q_reg_10 ( .CK(DNT_DW6_n126), .D(AD6IN_10), .R(TRST_), .Q(
        DW6[10]) );
    zdffqrb DNT_DW6_Q_reg_9 ( .CK(DNT_DW6_n126), .D(AD6IN_9), .R(TRST_), .Q(
        DW6[9]) );
    zdffqrb DNT_DW6_Q_reg_8 ( .CK(DNT_DW6_n126), .D(AD6IN_8), .R(TRST_), .Q(
        DW6[8]) );
    zdffqrb DNT_DW6_Q_reg_7 ( .CK(DNT_DW6_n126), .D(AD6IN_7), .R(TRST_), .Q(
        DW6[7]) );
    zdffqrb DNT_DW6_Q_reg_6 ( .CK(DNT_DW6_n126), .D(AD6IN_6), .R(TRST_), .Q(
        DW6[6]) );
    zdffqrb DNT_DW6_Q_reg_5 ( .CK(DNT_DW6_n126), .D(AD6IN_5), .R(TRST_), .Q(
        DW6[5]) );
    zdffqrb DNT_DW6_Q_reg_4 ( .CK(DNT_DW6_n126), .D(AD6IN_4), .R(TRST_), .Q(
        DW6[4]) );
    zdffqrb DNT_DW6_Q_reg_3 ( .CK(DNT_DW6_n126), .D(AD6IN_3), .R(TRST_), .Q(
        DW6[3]) );
    zdffqrb DNT_DW6_Q_reg_2 ( .CK(DNT_DW6_n126), .D(AD6IN_2), .R(TRST_), .Q(
        DW6[2]) );
    zdffqrb DNT_DW6_Q_reg_1 ( .CK(DNT_DW6_n126), .D(AD6IN_1), .R(TRST_), .Q(
        DW6[1]) );
    zdffqrb DNT_DW6_Q_reg_0 ( .CK(DNT_DW6_n126), .D(AD6IN_0), .R(TRST_), .Q(
        DW6[0]) );
    zbfb DNT_DW6_U80 ( .A(FLOPS_CLK_6), .Y(DNT_DW6_n126) );
    zbfb DNT_DW6_U81 ( .A(FLOPS_CLK_6), .Y(DNT_DW6_n127) );
    zdffqrb DNT_DW1_Q_reg_31 ( .CK(DNT_DW1_n127), .D(n445), .R(TRST_), .Q(DW1
        [31]) );
    zdffqrb DNT_DW1_Q_reg_30 ( .CK(DNT_DW1_n127), .D(n470), .R(TRST_), .Q(DW1
        [30]) );
    zdffqrb DNT_DW1_Q_reg_29 ( .CK(DNT_DW1_n127), .D(n475), .R(TRST_), .Q(DW1
        [29]) );
    zdffqrb DNT_DW1_Q_reg_28 ( .CK(DNT_DW1_n127), .D(n453), .R(TRST_), .Q(DW1
        [28]) );
    zdffqrb DNT_DW1_Q_reg_27 ( .CK(DNT_DW1_n127), .D(n465), .R(TRST_), .Q(DW1
        [27]) );
    zdffqrb DNT_DW1_Q_reg_26 ( .CK(DNT_DW1_n127), .D(n459), .R(TRST_), .Q(DW1
        [26]) );
    zdffqrb DNT_DW1_Q_reg_25 ( .CK(DNT_DW1_n127), .D(n464), .R(TRST_), .Q(DW1
        [25]) );
    zdffqrb DNT_DW1_Q_reg_24 ( .CK(DNT_DW1_n127), .D(n456), .R(TRST_), .Q(DW1
        [24]) );
    zdffqrb DNT_DW1_Q_reg_23 ( .CK(DNT_DW1_n127), .D(n449), .R(TRST_), .Q(DW1
        [23]) );
    zdffqrb DNT_DW1_Q_reg_22 ( .CK(DNT_DW1_n127), .D(n468), .R(TRST_), .Q(DW1
        [22]) );
    zdffqrb DNT_DW1_Q_reg_21 ( .CK(DNT_DW1_n127), .D(n457), .R(TRST_), .Q(DW1
        [21]) );
    zdffqrb DNT_DW1_Q_reg_20 ( .CK(DNT_DW1_n127), .D(n476), .R(TRST_), .Q(DW1
        [20]) );
    zdffqrb DNT_DW1_Q_reg_19 ( .CK(DNT_DW1_n127), .D(n466), .R(TRST_), .Q(DW1
        [19]) );
    zdffqrb DNT_DW1_Q_reg_18 ( .CK(DNT_DW1_n127), .D(n452), .R(TRST_), .Q(DW1
        [18]) );
    zdffqrb DNT_DW1_Q_reg_17 ( .CK(DNT_DW1_n127), .D(n472), .R(TRST_), .Q(DW1
        [17]) );
    zdffqrb DNT_DW1_Q_reg_16 ( .CK(DNT_DW1_n127), .D(n446), .R(TRST_), .Q(DW1
        [16]) );
    zdffqrb DNT_DW1_Q_reg_15 ( .CK(DNT_DW1_n126), .D(n471), .R(TRST_), .Q(DW1
        [15]) );
    zdffqrb DNT_DW1_Q_reg_14 ( .CK(DNT_DW1_n126), .D(n455), .R(TRST_), .Q(DW1
        [14]) );
    zdffqrb DNT_DW1_Q_reg_13 ( .CK(DNT_DW1_n126), .D(n461), .R(TRST_), .Q(DW1
        [13]) );
    zdffqrb DNT_DW1_Q_reg_12 ( .CK(DNT_DW1_n126), .D(n469), .R(TRST_), .Q(DW1
        [12]) );
    zdffqrb DNT_DW1_Q_reg_11 ( .CK(DNT_DW1_n126), .D(n448), .R(TRST_), .Q(DW1
        [11]) );
    zdffqrb DNT_DW1_Q_reg_10 ( .CK(DNT_DW1_n126), .D(n460), .R(TRST_), .Q(DW1
        [10]) );
    zdffqrb DNT_DW1_Q_reg_9 ( .CK(DNT_DW1_n126), .D(n454), .R(TRST_), .Q(DW1
        [9]) );
    zdffqrb DNT_DW1_Q_reg_8 ( .CK(DNT_DW1_n126), .D(n462), .R(TRST_), .Q(DW1
        [8]) );
    zdffqrb DNT_DW1_Q_reg_7 ( .CK(DNT_DW1_n126), .D(n447), .R(TRST_), .Q(DW1
        [7]) );
    zdffqrb DNT_DW1_Q_reg_6 ( .CK(DNT_DW1_n126), .D(n474), .R(TRST_), .Q(DW1
        [6]) );
    zdffqrb DNT_DW1_Q_reg_5 ( .CK(DNT_DW1_n126), .D(n451), .R(TRST_), .Q(DW1
        [5]) );
    zdffqrb DNT_DW1_Q_reg_4 ( .CK(DNT_DW1_n126), .D(n473), .R(TRST_), .Q(DW1
        [4]) );
    zdffqrb DNT_DW1_Q_reg_3 ( .CK(DNT_DW1_n126), .D(n467), .R(TRST_), .Q(DW1
        [3]) );
    zdffqrb DNT_DW1_Q_reg_2 ( .CK(DNT_DW1_n126), .D(n463), .R(TRST_), .Q(DW1
        [2]) );
    zdffqrb DNT_DW1_Q_reg_1 ( .CK(DNT_DW1_n126), .D(n458), .R(TRST_), .Q(DW1
        [1]) );
    zdffqrb DNT_DW1_Q_reg_0 ( .CK(DNT_DW1_n126), .D(n450), .R(TRST_), .Q(DW1
        [0]) );
    zbfb DNT_DW1_U80 ( .A(FLOPS_CLK_1), .Y(DNT_DW1_n126) );
    zbfb DNT_DW1_U81 ( .A(FLOPS_CLK_1), .Y(DNT_DW1_n127) );
    zdffqrb DNT_DW10_Q_reg_31 ( .CK(DNT_DW10_n127), .D(ADI[31]), .R(TRST_), 
        .Q(DW10[31]) );
    zdffqrb DNT_DW10_Q_reg_30 ( .CK(DNT_DW10_n127), .D(ADI[30]), .R(TRST_), 
        .Q(DW10[30]) );
    zdffqrb DNT_DW10_Q_reg_29 ( .CK(DNT_DW10_n127), .D(ADI[29]), .R(TRST_), 
        .Q(DW10[29]) );
    zdffqrb DNT_DW10_Q_reg_28 ( .CK(DNT_DW10_n127), .D(ADI[28]), .R(TRST_), 
        .Q(DW10[28]) );
    zdffqrb DNT_DW10_Q_reg_27 ( .CK(DNT_DW10_n127), .D(ADI[27]), .R(TRST_), 
        .Q(DW10[27]) );
    zdffqrb DNT_DW10_Q_reg_26 ( .CK(DNT_DW10_n127), .D(ADI[26]), .R(TRST_), 
        .Q(DW10[26]) );
    zdffqrb DNT_DW10_Q_reg_25 ( .CK(DNT_DW10_n127), .D(ADI[25]), .R(TRST_), 
        .Q(DW10[25]) );
    zdffqrb DNT_DW10_Q_reg_24 ( .CK(DNT_DW10_n127), .D(ADI[24]), .R(TRST_), 
        .Q(DW10[24]) );
    zdffqrb DNT_DW10_Q_reg_23 ( .CK(DNT_DW10_n127), .D(ADI[23]), .R(TRST_), 
        .Q(DW10[23]) );
    zdffqrb DNT_DW10_Q_reg_22 ( .CK(DNT_DW10_n127), .D(ADI[22]), .R(TRST_), 
        .Q(DW10[22]) );
    zdffqrb DNT_DW10_Q_reg_21 ( .CK(DNT_DW10_n127), .D(ADI[21]), .R(TRST_), 
        .Q(DW10[21]) );
    zdffqrb DNT_DW10_Q_reg_20 ( .CK(DNT_DW10_n127), .D(ADI[20]), .R(TRST_), 
        .Q(DW10[20]) );
    zdffqrb DNT_DW10_Q_reg_19 ( .CK(DNT_DW10_n127), .D(ADI[19]), .R(TRST_), 
        .Q(DW10[19]) );
    zdffqrb DNT_DW10_Q_reg_18 ( .CK(DNT_DW10_n127), .D(ADI[18]), .R(TRST_), 
        .Q(DW10[18]) );
    zdffqrb DNT_DW10_Q_reg_17 ( .CK(DNT_DW10_n127), .D(ADI[17]), .R(TRST_), 
        .Q(DW10[17]) );
    zdffqrb DNT_DW10_Q_reg_16 ( .CK(DNT_DW10_n127), .D(ADI[16]), .R(TRST_), 
        .Q(DW10[16]) );
    zdffqrb DNT_DW10_Q_reg_15 ( .CK(DNT_DW10_n126), .D(ADI[15]), .R(TRST_), 
        .Q(DW10[15]) );
    zdffqrb DNT_DW10_Q_reg_14 ( .CK(DNT_DW10_n126), .D(ADI[14]), .R(TRST_), 
        .Q(DW10[14]) );
    zdffqrb DNT_DW10_Q_reg_13 ( .CK(DNT_DW10_n126), .D(ADI[13]), .R(TRST_), 
        .Q(DW10[13]) );
    zdffqrb DNT_DW10_Q_reg_12 ( .CK(DNT_DW10_n126), .D(ADI[12]), .R(TRST_), 
        .Q(DW10[12]) );
    zdffqrb DNT_DW10_Q_reg_11 ( .CK(DNT_DW10_n126), .D(ADI[11]), .R(TRST_), 
        .Q(DW10[11]) );
    zdffqrb DNT_DW10_Q_reg_10 ( .CK(DNT_DW10_n126), .D(ADI[10]), .R(TRST_), 
        .Q(DW10[10]) );
    zdffqrb DNT_DW10_Q_reg_9 ( .CK(DNT_DW10_n126), .D(ADI[9]), .R(TRST_), .Q(
        DW10[9]) );
    zdffqrb DNT_DW10_Q_reg_8 ( .CK(DNT_DW10_n126), .D(ADI[8]), .R(TRST_), .Q(
        DW10[8]) );
    zdffqrb DNT_DW10_Q_reg_7 ( .CK(DNT_DW10_n126), .D(ADI[7]), .R(TRST_), .Q(
        DW10[7]) );
    zdffqrb DNT_DW10_Q_reg_6 ( .CK(DNT_DW10_n126), .D(ADI[6]), .R(TRST_), .Q(
        DW10[6]) );
    zdffqrb DNT_DW10_Q_reg_5 ( .CK(DNT_DW10_n126), .D(ADI[5]), .R(TRST_), .Q(
        DW10[5]) );
    zdffqrb DNT_DW10_Q_reg_4 ( .CK(DNT_DW10_n126), .D(ADI[4]), .R(TRST_), .Q(
        DW10[4]) );
    zdffqrb DNT_DW10_Q_reg_3 ( .CK(DNT_DW10_n126), .D(ADI[3]), .R(TRST_), .Q(
        DW10[3]) );
    zdffqrb DNT_DW10_Q_reg_2 ( .CK(DNT_DW10_n126), .D(ADI[2]), .R(TRST_), .Q(
        DW10[2]) );
    zdffqrb DNT_DW10_Q_reg_1 ( .CK(DNT_DW10_n126), .D(ADI[1]), .R(TRST_), .Q(
        DW10[1]) );
    zdffqrb DNT_DW10_Q_reg_0 ( .CK(DNT_DW10_n126), .D(ADI[0]), .R(TRST_), .Q(
        DW10[0]) );
    zbfb DNT_DW10_U80 ( .A(FLOPS_CLK_10), .Y(DNT_DW10_n126) );
    zbfb DNT_DW10_U81 ( .A(FLOPS_CLK_10), .Y(DNT_DW10_n127) );
    zdffqrb DNT_DW8_Q_reg_31 ( .CK(DNT_DW8_n127), .D(AD8IN_31), .R(TRST_), .Q(
        DW8[31]) );
    zdffqrb DNT_DW8_Q_reg_30 ( .CK(DNT_DW8_n127), .D(AD8IN_30), .R(TRST_), .Q(
        DW8[30]) );
    zdffqrb DNT_DW8_Q_reg_29 ( .CK(DNT_DW8_n127), .D(AD8IN_29), .R(TRST_), .Q(
        DW8[29]) );
    zdffqrb DNT_DW8_Q_reg_28 ( .CK(DNT_DW8_n127), .D(AD8IN_28), .R(TRST_), .Q(
        DW8[28]) );
    zdffqrb DNT_DW8_Q_reg_27 ( .CK(DNT_DW8_n127), .D(AD8IN_27), .R(TRST_), .Q(
        DW8[27]) );
    zdffqrb DNT_DW8_Q_reg_26 ( .CK(DNT_DW8_n127), .D(AD8IN_26), .R(TRST_), .Q(
        DW8[26]) );
    zdffqrb DNT_DW8_Q_reg_25 ( .CK(DNT_DW8_n127), .D(AD8IN_25), .R(TRST_), .Q(
        DW8[25]) );
    zdffqrb DNT_DW8_Q_reg_24 ( .CK(DNT_DW8_n127), .D(AD8IN_24), .R(TRST_), .Q(
        DW8[24]) );
    zdffqrb DNT_DW8_Q_reg_23 ( .CK(DNT_DW8_n127), .D(AD8IN_23), .R(TRST_), .Q(
        DW8[23]) );
    zdffqrb DNT_DW8_Q_reg_22 ( .CK(DNT_DW8_n127), .D(AD8IN_22), .R(TRST_), .Q(
        DW8[22]) );
    zdffqrb DNT_DW8_Q_reg_21 ( .CK(DNT_DW8_n127), .D(AD8IN_21), .R(TRST_), .Q(
        DW8[21]) );
    zdffqrb DNT_DW8_Q_reg_20 ( .CK(DNT_DW8_n127), .D(AD8IN_20), .R(TRST_), .Q(
        DW8[20]) );
    zdffqrb DNT_DW8_Q_reg_19 ( .CK(DNT_DW8_n127), .D(AD8IN_19), .R(TRST_), .Q(
        DW8[19]) );
    zdffqrb DNT_DW8_Q_reg_18 ( .CK(DNT_DW8_n127), .D(AD8IN_18), .R(TRST_), .Q(
        DW8[18]) );
    zdffqrb DNT_DW8_Q_reg_17 ( .CK(DNT_DW8_n127), .D(AD8IN_17), .R(TRST_), .Q(
        DW8[17]) );
    zdffqrb DNT_DW8_Q_reg_16 ( .CK(DNT_DW8_n127), .D(AD8IN_16), .R(TRST_), .Q(
        DW8[16]) );
    zdffqrb DNT_DW8_Q_reg_15 ( .CK(DNT_DW8_n126), .D(AD8IN_15), .R(TRST_), .Q(
        DW8[15]) );
    zdffqrb DNT_DW8_Q_reg_14 ( .CK(DNT_DW8_n126), .D(AD8IN_14), .R(TRST_), .Q(
        DW8[14]) );
    zdffqrb DNT_DW8_Q_reg_13 ( .CK(DNT_DW8_n126), .D(AD8IN_13), .R(TRST_), .Q(
        DW8[13]) );
    zdffqrb DNT_DW8_Q_reg_12 ( .CK(DNT_DW8_n126), .D(AD8IN_12), .R(TRST_), .Q(
        DW8[12]) );
    zdffqrb DNT_DW8_Q_reg_11 ( .CK(DNT_DW8_n126), .D(AD8IN_11), .R(TRST_), .Q(
        DW8[11]) );
    zdffqrb DNT_DW8_Q_reg_10 ( .CK(DNT_DW8_n126), .D(AD8IN_10), .R(TRST_), .Q(
        DW8[10]) );
    zdffqrb DNT_DW8_Q_reg_9 ( .CK(DNT_DW8_n126), .D(AD8IN_9), .R(TRST_), .Q(
        DW8[9]) );
    zdffqrb DNT_DW8_Q_reg_8 ( .CK(DNT_DW8_n126), .D(AD8IN_8), .R(TRST_), .Q(
        DW8[8]) );
    zdffqrb DNT_DW8_Q_reg_7 ( .CK(DNT_DW8_n126), .D(AD8IN_7), .R(TRST_), .Q(
        DW8[7]) );
    zdffqrb DNT_DW8_Q_reg_6 ( .CK(DNT_DW8_n126), .D(AD8IN_6), .R(TRST_), .Q(
        DW8[6]) );
    zdffqrb DNT_DW8_Q_reg_5 ( .CK(DNT_DW8_n126), .D(AD8IN_5), .R(TRST_), .Q(
        DW8[5]) );
    zdffqrb DNT_DW8_Q_reg_4 ( .CK(DNT_DW8_n126), .D(AD8IN_4), .R(TRST_), .Q(
        DW8[4]) );
    zdffqrb DNT_DW8_Q_reg_3 ( .CK(DNT_DW8_n126), .D(AD8IN_3), .R(TRST_), .Q(
        DW8[3]) );
    zdffqrb DNT_DW8_Q_reg_2 ( .CK(DNT_DW8_n126), .D(AD8IN_2), .R(TRST_), .Q(
        DW8[2]) );
    zdffqrb DNT_DW8_Q_reg_1 ( .CK(DNT_DW8_n126), .D(AD8IN_1), .R(TRST_), .Q(
        DW8[1]) );
    zdffqrb DNT_DW8_Q_reg_0 ( .CK(DNT_DW8_n126), .D(AD8IN_0), .R(TRST_), .Q(
        DW8[0]) );
    zbfb DNT_DW8_U80 ( .A(FLOPS_CLK_8), .Y(DNT_DW8_n126) );
    zbfb DNT_DW8_U81 ( .A(FLOPS_CLK_8), .Y(DNT_DW8_n127) );
    zdffqrb DNT_DW0_Q_reg_31 ( .CK(DNT_DW0_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW0[31]) );
    zdffqrb DNT_DW0_Q_reg_30 ( .CK(DNT_DW0_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW0[30]) );
    zdffqrb DNT_DW0_Q_reg_29 ( .CK(DNT_DW0_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW0[29]) );
    zdffqrb DNT_DW0_Q_reg_28 ( .CK(DNT_DW0_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW0[28]) );
    zdffqrb DNT_DW0_Q_reg_27 ( .CK(DNT_DW0_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW0[27]) );
    zdffqrb DNT_DW0_Q_reg_26 ( .CK(DNT_DW0_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW0[26]) );
    zdffqrb DNT_DW0_Q_reg_25 ( .CK(DNT_DW0_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW0[25]) );
    zdffqrb DNT_DW0_Q_reg_24 ( .CK(DNT_DW0_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW0[24]) );
    zdffqrb DNT_DW0_Q_reg_23 ( .CK(DNT_DW0_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW0[23]) );
    zdffqrb DNT_DW0_Q_reg_22 ( .CK(DNT_DW0_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW0[22]) );
    zdffqrb DNT_DW0_Q_reg_21 ( .CK(DNT_DW0_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW0[21]) );
    zdffqrb DNT_DW0_Q_reg_20 ( .CK(DNT_DW0_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW0[20]) );
    zdffqrb DNT_DW0_Q_reg_19 ( .CK(DNT_DW0_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW0[19]) );
    zdffqrb DNT_DW0_Q_reg_18 ( .CK(DNT_DW0_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW0[18]) );
    zdffqrb DNT_DW0_Q_reg_17 ( .CK(DNT_DW0_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW0[17]) );
    zdffqrb DNT_DW0_Q_reg_16 ( .CK(DNT_DW0_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW0[16]) );
    zdffqrb DNT_DW0_Q_reg_15 ( .CK(DNT_DW0_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW0[15]) );
    zdffqrb DNT_DW0_Q_reg_14 ( .CK(DNT_DW0_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW0[14]) );
    zdffqrb DNT_DW0_Q_reg_13 ( .CK(DNT_DW0_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW0[13]) );
    zdffqrb DNT_DW0_Q_reg_12 ( .CK(DNT_DW0_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW0[12]) );
    zdffqrb DNT_DW0_Q_reg_11 ( .CK(DNT_DW0_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW0[11]) );
    zdffqrb DNT_DW0_Q_reg_10 ( .CK(DNT_DW0_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW0[10]) );
    zdffqrb DNT_DW0_Q_reg_9 ( .CK(DNT_DW0_n126), .D(ADI[9]), .R(TRST_), .Q(DW0
        [9]) );
    zdffqrb DNT_DW0_Q_reg_8 ( .CK(DNT_DW0_n126), .D(ADI[8]), .R(TRST_), .Q(DW0
        [8]) );
    zdffqrb DNT_DW0_Q_reg_7 ( .CK(DNT_DW0_n126), .D(ADI[7]), .R(TRST_), .Q(DW0
        [7]) );
    zdffqrb DNT_DW0_Q_reg_6 ( .CK(DNT_DW0_n126), .D(ADI[6]), .R(TRST_), .Q(DW0
        [6]) );
    zdffqrb DNT_DW0_Q_reg_5 ( .CK(DNT_DW0_n126), .D(ADI[5]), .R(TRST_), .Q(DW0
        [5]) );
    zdffqrb DNT_DW0_Q_reg_4 ( .CK(DNT_DW0_n126), .D(ADI[4]), .R(TRST_), .Q(DW0
        [4]) );
    zdffqrb DNT_DW0_Q_reg_3 ( .CK(DNT_DW0_n126), .D(ADI[3]), .R(TRST_), .Q(DW0
        [3]) );
    zdffqrb DNT_DW0_Q_reg_2 ( .CK(DNT_DW0_n126), .D(ADI[2]), .R(TRST_), .Q(DW0
        [2]) );
    zdffqrb DNT_DW0_Q_reg_1 ( .CK(DNT_DW0_n126), .D(ADI[1]), .R(TRST_), .Q(DW0
        [1]) );
    zdffqrb DNT_DW0_Q_reg_0 ( .CK(DNT_DW0_n126), .D(ADI[0]), .R(TRST_), .Q(DW0
        [0]) );
    zbfb DNT_DW0_U80 ( .A(FLOPS_CLK_0), .Y(DNT_DW0_n126) );
    zbfb DNT_DW0_U81 ( .A(FLOPS_CLK_0), .Y(DNT_DW0_n127) );
    zdffqrb DNT_DW11_Q_reg_31 ( .CK(DNT_DW11_n127), .D(ADI[31]), .R(TRST_), 
        .Q(DW11[31]) );
    zdffqrb DNT_DW11_Q_reg_30 ( .CK(DNT_DW11_n127), .D(ADI[30]), .R(TRST_), 
        .Q(DW11[30]) );
    zdffqrb DNT_DW11_Q_reg_29 ( .CK(DNT_DW11_n127), .D(ADI[29]), .R(TRST_), 
        .Q(DW11[29]) );
    zdffqrb DNT_DW11_Q_reg_28 ( .CK(DNT_DW11_n127), .D(ADI[28]), .R(TRST_), 
        .Q(DW11[28]) );
    zdffqrb DNT_DW11_Q_reg_27 ( .CK(DNT_DW11_n127), .D(ADI[27]), .R(TRST_), 
        .Q(DW11[27]) );
    zdffqrb DNT_DW11_Q_reg_26 ( .CK(DNT_DW11_n127), .D(ADI[26]), .R(TRST_), 
        .Q(DW11[26]) );
    zdffqrb DNT_DW11_Q_reg_25 ( .CK(DNT_DW11_n127), .D(ADI[25]), .R(TRST_), 
        .Q(DW11[25]) );
    zdffqrb DNT_DW11_Q_reg_24 ( .CK(DNT_DW11_n127), .D(ADI[24]), .R(TRST_), 
        .Q(DW11[24]) );
    zdffqrb DNT_DW11_Q_reg_23 ( .CK(DNT_DW11_n127), .D(ADI[23]), .R(TRST_), 
        .Q(DW11[23]) );
    zdffqrb DNT_DW11_Q_reg_22 ( .CK(DNT_DW11_n127), .D(ADI[22]), .R(TRST_), 
        .Q(DW11[22]) );
    zdffqrb DNT_DW11_Q_reg_21 ( .CK(DNT_DW11_n127), .D(ADI[21]), .R(TRST_), 
        .Q(DW11[21]) );
    zdffqrb DNT_DW11_Q_reg_20 ( .CK(DNT_DW11_n127), .D(ADI[20]), .R(TRST_), 
        .Q(DW11[20]) );
    zdffqrb DNT_DW11_Q_reg_19 ( .CK(DNT_DW11_n127), .D(ADI[19]), .R(TRST_), 
        .Q(DW11[19]) );
    zdffqrb DNT_DW11_Q_reg_18 ( .CK(DNT_DW11_n127), .D(ADI[18]), .R(TRST_), 
        .Q(DW11[18]) );
    zdffqrb DNT_DW11_Q_reg_17 ( .CK(DNT_DW11_n127), .D(ADI[17]), .R(TRST_), 
        .Q(DW11[17]) );
    zdffqrb DNT_DW11_Q_reg_16 ( .CK(DNT_DW11_n127), .D(ADI[16]), .R(TRST_), 
        .Q(DW11[16]) );
    zdffqrb DNT_DW11_Q_reg_15 ( .CK(DNT_DW11_n126), .D(ADI[15]), .R(TRST_), 
        .Q(DW11[15]) );
    zdffqrb DNT_DW11_Q_reg_14 ( .CK(DNT_DW11_n126), .D(ADI[14]), .R(TRST_), 
        .Q(DW11[14]) );
    zdffqrb DNT_DW11_Q_reg_13 ( .CK(DNT_DW11_n126), .D(ADI[13]), .R(TRST_), 
        .Q(DW11[13]) );
    zdffqrb DNT_DW11_Q_reg_12 ( .CK(DNT_DW11_n126), .D(ADI[12]), .R(TRST_), 
        .Q(DW11[12]) );
    zdffqrb DNT_DW11_Q_reg_11 ( .CK(DNT_DW11_n126), .D(ADI[11]), .R(TRST_), 
        .Q(DW11[11]) );
    zdffqrb DNT_DW11_Q_reg_10 ( .CK(DNT_DW11_n126), .D(ADI[10]), .R(TRST_), 
        .Q(DW11[10]) );
    zdffqrb DNT_DW11_Q_reg_9 ( .CK(DNT_DW11_n126), .D(ADI[9]), .R(TRST_), .Q(
        DW11[9]) );
    zdffqrb DNT_DW11_Q_reg_8 ( .CK(DNT_DW11_n126), .D(ADI[8]), .R(TRST_), .Q(
        DW11[8]) );
    zdffqrb DNT_DW11_Q_reg_7 ( .CK(DNT_DW11_n126), .D(ADI[7]), .R(TRST_), .Q(
        DW11[7]) );
    zdffqrb DNT_DW11_Q_reg_6 ( .CK(DNT_DW11_n126), .D(ADI[6]), .R(TRST_), .Q(
        DW11[6]) );
    zdffqrb DNT_DW11_Q_reg_5 ( .CK(DNT_DW11_n126), .D(ADI[5]), .R(TRST_), .Q(
        DW11[5]) );
    zdffqrb DNT_DW11_Q_reg_4 ( .CK(DNT_DW11_n126), .D(ADI[4]), .R(TRST_), .Q(
        DW11[4]) );
    zdffqrb DNT_DW11_Q_reg_3 ( .CK(DNT_DW11_n126), .D(ADI[3]), .R(TRST_), .Q(
        DW11[3]) );
    zdffqrb DNT_DW11_Q_reg_2 ( .CK(DNT_DW11_n126), .D(ADI[2]), .R(TRST_), .Q(
        DW11[2]) );
    zdffqrb DNT_DW11_Q_reg_1 ( .CK(DNT_DW11_n126), .D(ADI[1]), .R(TRST_), .Q(
        DW11[1]) );
    zdffqrb DNT_DW11_Q_reg_0 ( .CK(DNT_DW11_n126), .D(ADI[0]), .R(TRST_), .Q(
        DW11[0]) );
    zbfb DNT_DW11_U80 ( .A(FLOPS_CLK_11), .Y(DNT_DW11_n126) );
    zbfb DNT_DW11_U81 ( .A(FLOPS_CLK_11), .Y(DNT_DW11_n127) );
    zdffqrb DNT_DW9_Q_reg_31 ( .CK(DNT_DW9_n127), .D(AD9IN_31), .R(TRST_), .Q(
        DW9[31]) );
    zdffqrb DNT_DW9_Q_reg_30 ( .CK(DNT_DW9_n127), .D(AD9IN_30), .R(TRST_), .Q(
        DW9[30]) );
    zdffqrb DNT_DW9_Q_reg_29 ( .CK(DNT_DW9_n127), .D(AD9IN_29), .R(TRST_), .Q(
        DW9[29]) );
    zdffqrb DNT_DW9_Q_reg_28 ( .CK(DNT_DW9_n127), .D(AD9IN_28), .R(TRST_), .Q(
        DW9[28]) );
    zdffqrb DNT_DW9_Q_reg_27 ( .CK(DNT_DW9_n127), .D(AD9IN_27), .R(TRST_), .Q(
        DW9[27]) );
    zdffqrb DNT_DW9_Q_reg_26 ( .CK(DNT_DW9_n127), .D(AD9IN_26), .R(TRST_), .Q(
        DW9[26]) );
    zdffqrb DNT_DW9_Q_reg_25 ( .CK(DNT_DW9_n127), .D(AD9IN_25), .R(TRST_), .Q(
        DW9[25]) );
    zdffqrb DNT_DW9_Q_reg_24 ( .CK(DNT_DW9_n127), .D(AD9IN_24), .R(TRST_), .Q(
        DW9[24]) );
    zdffqrb DNT_DW9_Q_reg_23 ( .CK(DNT_DW9_n127), .D(AD9IN_23), .R(TRST_), .Q(
        DW9[23]) );
    zdffqrb DNT_DW9_Q_reg_22 ( .CK(DNT_DW9_n127), .D(AD9IN_22), .R(TRST_), .Q(
        DW9[22]) );
    zdffqrb DNT_DW9_Q_reg_21 ( .CK(DNT_DW9_n127), .D(AD9IN_21), .R(TRST_), .Q(
        DW9[21]) );
    zdffqrb DNT_DW9_Q_reg_20 ( .CK(DNT_DW9_n127), .D(AD9IN_20), .R(TRST_), .Q(
        DW9[20]) );
    zdffqrb DNT_DW9_Q_reg_19 ( .CK(DNT_DW9_n127), .D(AD9IN_19), .R(TRST_), .Q(
        DW9[19]) );
    zdffqrb DNT_DW9_Q_reg_18 ( .CK(DNT_DW9_n127), .D(AD9IN_18), .R(TRST_), .Q(
        DW9[18]) );
    zdffqrb DNT_DW9_Q_reg_17 ( .CK(DNT_DW9_n127), .D(AD9IN_17), .R(TRST_), .Q(
        DW9[17]) );
    zdffqrb DNT_DW9_Q_reg_16 ( .CK(DNT_DW9_n127), .D(AD9IN_16), .R(TRST_), .Q(
        DW9[16]) );
    zdffqrb DNT_DW9_Q_reg_15 ( .CK(DNT_DW9_n126), .D(AD9IN_15), .R(TRST_), .Q(
        DW9[15]) );
    zdffqrb DNT_DW9_Q_reg_14 ( .CK(DNT_DW9_n126), .D(AD9IN_14), .R(TRST_), .Q(
        DW9[14]) );
    zdffqrb DNT_DW9_Q_reg_13 ( .CK(DNT_DW9_n126), .D(AD9IN_13), .R(TRST_), .Q(
        DW9[13]) );
    zdffqrb DNT_DW9_Q_reg_12 ( .CK(DNT_DW9_n126), .D(AD9IN_12), .R(TRST_), .Q(
        DW9[12]) );
    zdffqrb DNT_DW9_Q_reg_11 ( .CK(DNT_DW9_n126), .D(AD9IN_11), .R(TRST_), .Q(
        DW9[11]) );
    zdffqrb DNT_DW9_Q_reg_10 ( .CK(DNT_DW9_n126), .D(AD9IN_10), .R(TRST_), .Q(
        DW9[10]) );
    zdffqrb DNT_DW9_Q_reg_9 ( .CK(DNT_DW9_n126), .D(AD9IN_9), .R(TRST_), .Q(
        DW9[9]) );
    zdffqrb DNT_DW9_Q_reg_8 ( .CK(DNT_DW9_n126), .D(AD9IN_8), .R(TRST_), .Q(
        DW9[8]) );
    zdffqrb DNT_DW9_Q_reg_7 ( .CK(DNT_DW9_n126), .D(AD9IN_7), .R(TRST_), .Q(
        DW9[7]) );
    zdffqrb DNT_DW9_Q_reg_6 ( .CK(DNT_DW9_n126), .D(AD9IN_6), .R(TRST_), .Q(
        DW9[6]) );
    zdffqrb DNT_DW9_Q_reg_5 ( .CK(DNT_DW9_n126), .D(AD9IN_5), .R(TRST_), .Q(
        DW9[5]) );
    zdffqrb DNT_DW9_Q_reg_4 ( .CK(DNT_DW9_n126), .D(AD9IN_4), .R(TRST_), .Q(
        DW9[4]) );
    zdffqrb DNT_DW9_Q_reg_3 ( .CK(DNT_DW9_n126), .D(AD9IN_3), .R(TRST_), .Q(
        DW9[3]) );
    zdffqrb DNT_DW9_Q_reg_2 ( .CK(DNT_DW9_n126), .D(AD9IN_2), .R(TRST_), .Q(
        DW9[2]) );
    zdffqrb DNT_DW9_Q_reg_1 ( .CK(DNT_DW9_n126), .D(AD9IN_1), .R(TRST_), .Q(
        DW9[1]) );
    zdffqrb DNT_DW9_Q_reg_0 ( .CK(DNT_DW9_n126), .D(AD9IN_0), .R(TRST_), .Q(
        DW9[0]) );
    zbfb DNT_DW9_U80 ( .A(FLOPS_CLK_9), .Y(DNT_DW9_n126) );
    zbfb DNT_DW9_U81 ( .A(FLOPS_CLK_9), .Y(DNT_DW9_n127) );
    zdffqrb DNT_DW7_Q_reg_31 ( .CK(DNT_DW7_n127), .D(AD7IN_31), .R(TRST_), .Q(
        DW7[31]) );
    zdffqrb DNT_DW7_Q_reg_30 ( .CK(DNT_DW7_n127), .D(AD7IN_30), .R(TRST_), .Q(
        DW7[30]) );
    zdffqrb DNT_DW7_Q_reg_29 ( .CK(DNT_DW7_n127), .D(AD7IN_29), .R(TRST_), .Q(
        DW7[29]) );
    zdffqrb DNT_DW7_Q_reg_28 ( .CK(DNT_DW7_n127), .D(AD7IN_28), .R(TRST_), .Q(
        DW7[28]) );
    zdffqrb DNT_DW7_Q_reg_27 ( .CK(DNT_DW7_n127), .D(AD7IN_27), .R(TRST_), .Q(
        DW7[27]) );
    zdffqrb DNT_DW7_Q_reg_26 ( .CK(DNT_DW7_n127), .D(AD7IN_26), .R(TRST_), .Q(
        DW7[26]) );
    zdffqrb DNT_DW7_Q_reg_25 ( .CK(DNT_DW7_n127), .D(AD7IN_25), .R(TRST_), .Q(
        DW7[25]) );
    zdffqrb DNT_DW7_Q_reg_24 ( .CK(DNT_DW7_n127), .D(AD7IN_24), .R(TRST_), .Q(
        DW7[24]) );
    zdffqrb DNT_DW7_Q_reg_23 ( .CK(DNT_DW7_n127), .D(AD7IN_23), .R(TRST_), .Q(
        DW7[23]) );
    zdffqrb DNT_DW7_Q_reg_22 ( .CK(DNT_DW7_n127), .D(AD7IN_22), .R(TRST_), .Q(
        DW7[22]) );
    zdffqrb DNT_DW7_Q_reg_21 ( .CK(DNT_DW7_n127), .D(AD7IN_21), .R(TRST_), .Q(
        DW7[21]) );
    zdffqrb DNT_DW7_Q_reg_20 ( .CK(DNT_DW7_n127), .D(AD7IN_20), .R(TRST_), .Q(
        DW7[20]) );
    zdffqrb DNT_DW7_Q_reg_19 ( .CK(DNT_DW7_n127), .D(AD7IN_19), .R(TRST_), .Q(
        DW7[19]) );
    zdffqrb DNT_DW7_Q_reg_18 ( .CK(DNT_DW7_n127), .D(AD7IN_18), .R(TRST_), .Q(
        DW7[18]) );
    zdffqrb DNT_DW7_Q_reg_17 ( .CK(DNT_DW7_n127), .D(AD7IN_17), .R(TRST_), .Q(
        DW7[17]) );
    zdffqrb DNT_DW7_Q_reg_16 ( .CK(DNT_DW7_n127), .D(AD7IN_16), .R(TRST_), .Q(
        DW7[16]) );
    zdffqrb DNT_DW7_Q_reg_15 ( .CK(DNT_DW7_n126), .D(AD7IN_15), .R(TRST_), .Q(
        DW7[15]) );
    zdffqrb DNT_DW7_Q_reg_14 ( .CK(DNT_DW7_n126), .D(AD7IN_14), .R(TRST_), .Q(
        DW7[14]) );
    zdffqrb DNT_DW7_Q_reg_13 ( .CK(DNT_DW7_n126), .D(AD7IN_13), .R(TRST_), .Q(
        DW7[13]) );
    zdffqrb DNT_DW7_Q_reg_12 ( .CK(DNT_DW7_n126), .D(AD7IN_12), .R(TRST_), .Q(
        DW7[12]) );
    zdffqrb DNT_DW7_Q_reg_11 ( .CK(DNT_DW7_n126), .D(AD7IN_11), .R(TRST_), .Q(
        DW7[11]) );
    zdffqrb DNT_DW7_Q_reg_10 ( .CK(DNT_DW7_n126), .D(AD7IN_10), .R(TRST_), .Q(
        DW7[10]) );
    zdffqrb DNT_DW7_Q_reg_9 ( .CK(DNT_DW7_n126), .D(AD7IN_9), .R(TRST_), .Q(
        DW7[9]) );
    zdffqrb DNT_DW7_Q_reg_8 ( .CK(DNT_DW7_n126), .D(AD7IN_8), .R(TRST_), .Q(
        DW7[8]) );
    zdffqrb DNT_DW7_Q_reg_7 ( .CK(DNT_DW7_n126), .D(AD7IN_7), .R(TRST_), .Q(
        DW7[7]) );
    zdffqrb DNT_DW7_Q_reg_6 ( .CK(DNT_DW7_n126), .D(AD7IN_6), .R(TRST_), .Q(
        DW7[6]) );
    zdffqrb DNT_DW7_Q_reg_5 ( .CK(DNT_DW7_n126), .D(AD7IN_5), .R(TRST_), .Q(
        DW7[5]) );
    zdffqrb DNT_DW7_Q_reg_4 ( .CK(DNT_DW7_n126), .D(AD7IN_4), .R(TRST_), .Q(
        DW7[4]) );
    zdffqrb DNT_DW7_Q_reg_3 ( .CK(DNT_DW7_n126), .D(AD7IN_3), .R(TRST_), .Q(
        DW7[3]) );
    zdffqrb DNT_DW7_Q_reg_2 ( .CK(DNT_DW7_n126), .D(AD7IN_2), .R(TRST_), .Q(
        DW7[2]) );
    zdffqrb DNT_DW7_Q_reg_1 ( .CK(DNT_DW7_n126), .D(AD7IN_1), .R(TRST_), .Q(
        DW7[1]) );
    zdffqrb DNT_DW7_Q_reg_0 ( .CK(DNT_DW7_n126), .D(AD7IN_0), .R(TRST_), .Q(
        DW7[0]) );
    zbfb DNT_DW7_U80 ( .A(FLOPS_CLK_7), .Y(DNT_DW7_n126) );
    zbfb DNT_DW7_U81 ( .A(FLOPS_CLK_7), .Y(DNT_DW7_n127) );
    zdffqrb DNT_DW5_Q_reg_31 ( .CK(DNT_DW5_n127), .D(AD5IN_31), .R(TRST_), .Q(
        DW5[31]) );
    zdffqrb DNT_DW5_Q_reg_30 ( .CK(DNT_DW5_n127), .D(AD5IN_30), .R(TRST_), .Q(
        DW5[30]) );
    zdffqrb DNT_DW5_Q_reg_29 ( .CK(DNT_DW5_n127), .D(AD5IN_29), .R(TRST_), .Q(
        DW5[29]) );
    zdffqrb DNT_DW5_Q_reg_28 ( .CK(DNT_DW5_n127), .D(AD5IN_28), .R(TRST_), .Q(
        DW5[28]) );
    zdffqrb DNT_DW5_Q_reg_27 ( .CK(DNT_DW5_n127), .D(AD5IN_27), .R(TRST_), .Q(
        DW5[27]) );
    zdffqrb DNT_DW5_Q_reg_26 ( .CK(DNT_DW5_n127), .D(AD5IN_26), .R(TRST_), .Q(
        DW5[26]) );
    zdffqrb DNT_DW5_Q_reg_25 ( .CK(DNT_DW5_n127), .D(AD5IN_25), .R(TRST_), .Q(
        DW5[25]) );
    zdffqrb DNT_DW5_Q_reg_24 ( .CK(DNT_DW5_n127), .D(AD5IN_24), .R(TRST_), .Q(
        DW5[24]) );
    zdffqrb DNT_DW5_Q_reg_23 ( .CK(DNT_DW5_n127), .D(AD5IN_23), .R(TRST_), .Q(
        DW5[23]) );
    zdffqrb DNT_DW5_Q_reg_22 ( .CK(DNT_DW5_n127), .D(AD5IN_22), .R(TRST_), .Q(
        DW5[22]) );
    zdffqrb DNT_DW5_Q_reg_21 ( .CK(DNT_DW5_n127), .D(AD5IN_21), .R(TRST_), .Q(
        DW5[21]) );
    zdffqrb DNT_DW5_Q_reg_20 ( .CK(DNT_DW5_n127), .D(AD5IN_20), .R(TRST_), .Q(
        DW5[20]) );
    zdffqrb DNT_DW5_Q_reg_19 ( .CK(DNT_DW5_n127), .D(AD5IN_19), .R(TRST_), .Q(
        DW5[19]) );
    zdffqrb DNT_DW5_Q_reg_18 ( .CK(DNT_DW5_n127), .D(AD5IN_18), .R(TRST_), .Q(
        DW5[18]) );
    zdffqrb DNT_DW5_Q_reg_17 ( .CK(DNT_DW5_n127), .D(AD5IN_17), .R(TRST_), .Q(
        DW5[17]) );
    zdffqrb DNT_DW5_Q_reg_16 ( .CK(DNT_DW5_n127), .D(AD5IN_16), .R(TRST_), .Q(
        DW5[16]) );
    zdffqrb DNT_DW5_Q_reg_15 ( .CK(DNT_DW5_n126), .D(AD5IN_15), .R(TRST_), .Q(
        DW5[15]) );
    zdffqrb DNT_DW5_Q_reg_14 ( .CK(DNT_DW5_n126), .D(AD5IN_14), .R(TRST_), .Q(
        DW5[14]) );
    zdffqrb DNT_DW5_Q_reg_13 ( .CK(DNT_DW5_n126), .D(AD5IN_13), .R(TRST_), .Q(
        DW5[13]) );
    zdffqrb DNT_DW5_Q_reg_12 ( .CK(DNT_DW5_n126), .D(AD5IN_12), .R(TRST_), .Q(
        DW5[12]) );
    zdffqrb DNT_DW5_Q_reg_11 ( .CK(DNT_DW5_n126), .D(AD5IN_11), .R(TRST_), .Q(
        DW5[11]) );
    zdffqrb DNT_DW5_Q_reg_10 ( .CK(DNT_DW5_n126), .D(AD5IN_10), .R(TRST_), .Q(
        DW5[10]) );
    zdffqrb DNT_DW5_Q_reg_9 ( .CK(DNT_DW5_n126), .D(AD5IN_9), .R(TRST_), .Q(
        DW5[9]) );
    zdffqrb DNT_DW5_Q_reg_8 ( .CK(DNT_DW5_n126), .D(AD5IN_8), .R(TRST_), .Q(
        DW5[8]) );
    zdffqrb DNT_DW5_Q_reg_7 ( .CK(DNT_DW5_n126), .D(AD5IN_7), .R(TRST_), .Q(
        DW5[7]) );
    zdffqrb DNT_DW5_Q_reg_6 ( .CK(DNT_DW5_n126), .D(AD5IN_6), .R(TRST_), .Q(
        DW5[6]) );
    zdffqrb DNT_DW5_Q_reg_5 ( .CK(DNT_DW5_n126), .D(AD5IN_5), .R(TRST_), .Q(
        DW5[5]) );
    zdffqrb DNT_DW5_Q_reg_4 ( .CK(DNT_DW5_n126), .D(AD5IN_4), .R(TRST_), .Q(
        DW5[4]) );
    zdffqrb DNT_DW5_Q_reg_3 ( .CK(DNT_DW5_n126), .D(AD5IN_3), .R(TRST_), .Q(
        DW5[3]) );
    zdffqrb DNT_DW5_Q_reg_2 ( .CK(DNT_DW5_n126), .D(AD5IN_2), .R(TRST_), .Q(
        DW5[2]) );
    zdffqrb DNT_DW5_Q_reg_1 ( .CK(DNT_DW5_n126), .D(AD5IN_1), .R(TRST_), .Q(
        DW5[1]) );
    zdffqrb DNT_DW5_Q_reg_0 ( .CK(DNT_DW5_n126), .D(AD5IN_0), .R(TRST_), .Q(
        DW5[0]) );
    zbfb DNT_DW5_U80 ( .A(FLOPS_CLK_5), .Y(DNT_DW5_n126) );
    zbfb DNT_DW5_U81 ( .A(FLOPS_CLK_5), .Y(DNT_DW5_n127) );
    zdffqrb DNT_DW14_Q_reg_31 ( .CK(DNT_DW14_n127), .D(ADI[31]), .R(TRST_), 
        .Q(DW14[31]) );
    zdffqrb DNT_DW14_Q_reg_30 ( .CK(DNT_DW14_n127), .D(ADI[30]), .R(TRST_), 
        .Q(DW14[30]) );
    zdffqrb DNT_DW14_Q_reg_29 ( .CK(DNT_DW14_n127), .D(ADI[29]), .R(TRST_), 
        .Q(DW14[29]) );
    zdffqrb DNT_DW14_Q_reg_28 ( .CK(DNT_DW14_n127), .D(ADI[28]), .R(TRST_), 
        .Q(DW14[28]) );
    zdffqrb DNT_DW14_Q_reg_27 ( .CK(DNT_DW14_n127), .D(ADI[27]), .R(TRST_), 
        .Q(DW14[27]) );
    zdffqrb DNT_DW14_Q_reg_26 ( .CK(DNT_DW14_n127), .D(ADI[26]), .R(TRST_), 
        .Q(DW14[26]) );
    zdffqrb DNT_DW14_Q_reg_25 ( .CK(DNT_DW14_n127), .D(ADI[25]), .R(TRST_), 
        .Q(DW14[25]) );
    zdffqrb DNT_DW14_Q_reg_24 ( .CK(DNT_DW14_n127), .D(ADI[24]), .R(TRST_), 
        .Q(DW14[24]) );
    zdffqrb DNT_DW14_Q_reg_23 ( .CK(DNT_DW14_n127), .D(ADI[23]), .R(TRST_), 
        .Q(DW14[23]) );
    zdffqrb DNT_DW14_Q_reg_22 ( .CK(DNT_DW14_n127), .D(ADI[22]), .R(TRST_), 
        .Q(DW14[22]) );
    zdffqrb DNT_DW14_Q_reg_21 ( .CK(DNT_DW14_n127), .D(ADI[21]), .R(TRST_), 
        .Q(DW14[21]) );
    zdffqrb DNT_DW14_Q_reg_20 ( .CK(DNT_DW14_n127), .D(ADI[20]), .R(TRST_), 
        .Q(DW14[20]) );
    zdffqrb DNT_DW14_Q_reg_19 ( .CK(DNT_DW14_n127), .D(ADI[19]), .R(TRST_), 
        .Q(DW14[19]) );
    zdffqrb DNT_DW14_Q_reg_18 ( .CK(DNT_DW14_n127), .D(ADI[18]), .R(TRST_), 
        .Q(DW14[18]) );
    zdffqrb DNT_DW14_Q_reg_17 ( .CK(DNT_DW14_n127), .D(ADI[17]), .R(TRST_), 
        .Q(DW14[17]) );
    zdffqrb DNT_DW14_Q_reg_16 ( .CK(DNT_DW14_n127), .D(ADI[16]), .R(TRST_), 
        .Q(DW14[16]) );
    zdffqrb DNT_DW14_Q_reg_15 ( .CK(DNT_DW14_n126), .D(ADI[15]), .R(TRST_), 
        .Q(DW14[15]) );
    zdffqrb DNT_DW14_Q_reg_14 ( .CK(DNT_DW14_n126), .D(ADI[14]), .R(TRST_), 
        .Q(DW14[14]) );
    zdffqrb DNT_DW14_Q_reg_13 ( .CK(DNT_DW14_n126), .D(ADI[13]), .R(TRST_), 
        .Q(DW14[13]) );
    zdffqrb DNT_DW14_Q_reg_12 ( .CK(DNT_DW14_n126), .D(ADI[12]), .R(TRST_), 
        .Q(DW14[12]) );
    zdffqrb DNT_DW14_Q_reg_11 ( .CK(DNT_DW14_n126), .D(ADI[11]), .R(TRST_), 
        .Q(DW14[11]) );
    zdffqrb DNT_DW14_Q_reg_10 ( .CK(DNT_DW14_n126), .D(ADI[10]), .R(TRST_), 
        .Q(DW14[10]) );
    zdffqrb DNT_DW14_Q_reg_9 ( .CK(DNT_DW14_n126), .D(ADI[9]), .R(TRST_), .Q(
        DW14[9]) );
    zdffqrb DNT_DW14_Q_reg_8 ( .CK(DNT_DW14_n126), .D(ADI[8]), .R(TRST_), .Q(
        DW14[8]) );
    zdffqrb DNT_DW14_Q_reg_7 ( .CK(DNT_DW14_n126), .D(ADI[7]), .R(TRST_), .Q(
        DW14[7]) );
    zdffqrb DNT_DW14_Q_reg_6 ( .CK(DNT_DW14_n126), .D(ADI[6]), .R(TRST_), .Q(
        DW14[6]) );
    zdffqrb DNT_DW14_Q_reg_5 ( .CK(DNT_DW14_n126), .D(ADI[5]), .R(TRST_), .Q(
        DW14[5]) );
    zdffqrb DNT_DW14_Q_reg_4 ( .CK(DNT_DW14_n126), .D(ADI[4]), .R(TRST_), .Q(
        DW14[4]) );
    zdffqrb DNT_DW14_Q_reg_3 ( .CK(DNT_DW14_n126), .D(ADI[3]), .R(TRST_), .Q(
        DW14[3]) );
    zdffqrb DNT_DW14_Q_reg_2 ( .CK(DNT_DW14_n126), .D(ADI[2]), .R(TRST_), .Q(
        DW14[2]) );
    zdffqrb DNT_DW14_Q_reg_1 ( .CK(DNT_DW14_n126), .D(ADI[1]), .R(TRST_), .Q(
        DW14[1]) );
    zdffqrb DNT_DW14_Q_reg_0 ( .CK(DNT_DW14_n126), .D(ADI[0]), .R(TRST_), .Q(
        DW14[0]) );
    zbfb DNT_DW14_U80 ( .A(FLOPS_CLK_14), .Y(DNT_DW14_n126) );
    zbfb DNT_DW14_U81 ( .A(FLOPS_CLK_14), .Y(DNT_DW14_n127) );
    zdffqrb DNT_DW2_Q_reg_31 ( .CK(DNT_DW2_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW2[31]) );
    zdffqrb DNT_DW2_Q_reg_30 ( .CK(DNT_DW2_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW2[30]) );
    zdffqrb DNT_DW2_Q_reg_29 ( .CK(DNT_DW2_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW2[29]) );
    zdffqrb DNT_DW2_Q_reg_28 ( .CK(DNT_DW2_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW2[28]) );
    zdffqrb DNT_DW2_Q_reg_27 ( .CK(DNT_DW2_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW2[27]) );
    zdffqrb DNT_DW2_Q_reg_26 ( .CK(DNT_DW2_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW2[26]) );
    zdffqrb DNT_DW2_Q_reg_25 ( .CK(DNT_DW2_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW2[25]) );
    zdffqrb DNT_DW2_Q_reg_24 ( .CK(DNT_DW2_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW2[24]) );
    zdffqrb DNT_DW2_Q_reg_23 ( .CK(DNT_DW2_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW2[23]) );
    zdffqrb DNT_DW2_Q_reg_22 ( .CK(DNT_DW2_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW2[22]) );
    zdffqrb DNT_DW2_Q_reg_21 ( .CK(DNT_DW2_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW2[21]) );
    zdffqrb DNT_DW2_Q_reg_20 ( .CK(DNT_DW2_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW2[20]) );
    zdffqrb DNT_DW2_Q_reg_19 ( .CK(DNT_DW2_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW2[19]) );
    zdffqrb DNT_DW2_Q_reg_18 ( .CK(DNT_DW2_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW2[18]) );
    zdffqrb DNT_DW2_Q_reg_17 ( .CK(DNT_DW2_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW2[17]) );
    zdffqrb DNT_DW2_Q_reg_16 ( .CK(DNT_DW2_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW2[16]) );
    zdffqrb DNT_DW2_Q_reg_15 ( .CK(DNT_DW2_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW2[15]) );
    zdffqrb DNT_DW2_Q_reg_14 ( .CK(DNT_DW2_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW2[14]) );
    zdffqrb DNT_DW2_Q_reg_13 ( .CK(DNT_DW2_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW2[13]) );
    zdffqrb DNT_DW2_Q_reg_12 ( .CK(DNT_DW2_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW2[12]) );
    zdffqrb DNT_DW2_Q_reg_11 ( .CK(DNT_DW2_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW2[11]) );
    zdffqrb DNT_DW2_Q_reg_10 ( .CK(DNT_DW2_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW2[10]) );
    zdffqrb DNT_DW2_Q_reg_9 ( .CK(DNT_DW2_n126), .D(ADI[9]), .R(TRST_), .Q(DW2
        [9]) );
    zdffqrb DNT_DW2_Q_reg_8 ( .CK(DNT_DW2_n126), .D(ADI[8]), .R(TRST_), .Q(DW2
        [8]) );
    zdffqrb DNT_DW2_Q_reg_7 ( .CK(DNT_DW2_n126), .D(ADI[7]), .R(TRST_), .Q(DW2
        [7]) );
    zdffqrb DNT_DW2_Q_reg_6 ( .CK(DNT_DW2_n126), .D(ADI[6]), .R(TRST_), .Q(DW2
        [6]) );
    zdffqrb DNT_DW2_Q_reg_5 ( .CK(DNT_DW2_n126), .D(ADI[5]), .R(TRST_), .Q(DW2
        [5]) );
    zdffqrb DNT_DW2_Q_reg_4 ( .CK(DNT_DW2_n126), .D(ADI[4]), .R(TRST_), .Q(DW2
        [4]) );
    zdffqrb DNT_DW2_Q_reg_3 ( .CK(DNT_DW2_n126), .D(ADI[3]), .R(TRST_), .Q(DW2
        [3]) );
    zdffqrb DNT_DW2_Q_reg_2 ( .CK(DNT_DW2_n126), .D(ADI[2]), .R(TRST_), .Q(DW2
        [2]) );
    zdffqrb DNT_DW2_Q_reg_1 ( .CK(DNT_DW2_n126), .D(ADI[1]), .R(TRST_), .Q(DW2
        [1]) );
    zdffqrb DNT_DW2_Q_reg_0 ( .CK(DNT_DW2_n126), .D(ADI[0]), .R(TRST_), .Q(DW2
        [0]) );
    zbfb DNT_DW2_U80 ( .A(FLOPS_CLK_2), .Y(DNT_DW2_n126) );
    zbfb DNT_DW2_U81 ( .A(FLOPS_CLK_2), .Y(DNT_DW2_n127) );
    zdffqrb DNT_DW13_Q_reg_31 ( .CK(DNT_DW13_n127), .D(ADI[31]), .R(TRST_), 
        .Q(DW13[31]) );
    zdffqrb DNT_DW13_Q_reg_30 ( .CK(DNT_DW13_n127), .D(ADI[30]), .R(TRST_), 
        .Q(DW13[30]) );
    zdffqrb DNT_DW13_Q_reg_29 ( .CK(DNT_DW13_n127), .D(ADI[29]), .R(TRST_), 
        .Q(DW13[29]) );
    zdffqrb DNT_DW13_Q_reg_28 ( .CK(DNT_DW13_n127), .D(ADI[28]), .R(TRST_), 
        .Q(DW13[28]) );
    zdffqrb DNT_DW13_Q_reg_27 ( .CK(DNT_DW13_n127), .D(ADI[27]), .R(TRST_), 
        .Q(DW13[27]) );
    zdffqrb DNT_DW13_Q_reg_26 ( .CK(DNT_DW13_n127), .D(ADI[26]), .R(TRST_), 
        .Q(DW13[26]) );
    zdffqrb DNT_DW13_Q_reg_25 ( .CK(DNT_DW13_n127), .D(ADI[25]), .R(TRST_), 
        .Q(DW13[25]) );
    zdffqrb DNT_DW13_Q_reg_24 ( .CK(DNT_DW13_n127), .D(ADI[24]), .R(TRST_), 
        .Q(DW13[24]) );
    zdffqrb DNT_DW13_Q_reg_23 ( .CK(DNT_DW13_n127), .D(ADI[23]), .R(TRST_), 
        .Q(DW13[23]) );
    zdffqrb DNT_DW13_Q_reg_22 ( .CK(DNT_DW13_n127), .D(ADI[22]), .R(TRST_), 
        .Q(DW13[22]) );
    zdffqrb DNT_DW13_Q_reg_21 ( .CK(DNT_DW13_n127), .D(ADI[21]), .R(TRST_), 
        .Q(DW13[21]) );
    zdffqrb DNT_DW13_Q_reg_20 ( .CK(DNT_DW13_n127), .D(ADI[20]), .R(TRST_), 
        .Q(DW13[20]) );
    zdffqrb DNT_DW13_Q_reg_19 ( .CK(DNT_DW13_n127), .D(ADI[19]), .R(TRST_), 
        .Q(DW13[19]) );
    zdffqrb DNT_DW13_Q_reg_18 ( .CK(DNT_DW13_n127), .D(ADI[18]), .R(TRST_), 
        .Q(DW13[18]) );
    zdffqrb DNT_DW13_Q_reg_17 ( .CK(DNT_DW13_n127), .D(ADI[17]), .R(TRST_), 
        .Q(DW13[17]) );
    zdffqrb DNT_DW13_Q_reg_16 ( .CK(DNT_DW13_n127), .D(ADI[16]), .R(TRST_), 
        .Q(DW13[16]) );
    zdffqrb DNT_DW13_Q_reg_15 ( .CK(DNT_DW13_n126), .D(ADI[15]), .R(TRST_), 
        .Q(DW13[15]) );
    zdffqrb DNT_DW13_Q_reg_14 ( .CK(DNT_DW13_n126), .D(ADI[14]), .R(TRST_), 
        .Q(DW13[14]) );
    zdffqrb DNT_DW13_Q_reg_13 ( .CK(DNT_DW13_n126), .D(ADI[13]), .R(TRST_), 
        .Q(DW13[13]) );
    zdffqrb DNT_DW13_Q_reg_12 ( .CK(DNT_DW13_n126), .D(ADI[12]), .R(TRST_), 
        .Q(DW13[12]) );
    zdffqrb DNT_DW13_Q_reg_11 ( .CK(DNT_DW13_n126), .D(ADI[11]), .R(TRST_), 
        .Q(DW13[11]) );
    zdffqrb DNT_DW13_Q_reg_10 ( .CK(DNT_DW13_n126), .D(ADI[10]), .R(TRST_), 
        .Q(DW13[10]) );
    zdffqrb DNT_DW13_Q_reg_9 ( .CK(DNT_DW13_n126), .D(ADI[9]), .R(TRST_), .Q(
        DW13[9]) );
    zdffqrb DNT_DW13_Q_reg_8 ( .CK(DNT_DW13_n126), .D(ADI[8]), .R(TRST_), .Q(
        DW13[8]) );
    zdffqrb DNT_DW13_Q_reg_7 ( .CK(DNT_DW13_n126), .D(ADI[7]), .R(TRST_), .Q(
        DW13[7]) );
    zdffqrb DNT_DW13_Q_reg_6 ( .CK(DNT_DW13_n126), .D(ADI[6]), .R(TRST_), .Q(
        DW13[6]) );
    zdffqrb DNT_DW13_Q_reg_5 ( .CK(DNT_DW13_n126), .D(ADI[5]), .R(TRST_), .Q(
        DW13[5]) );
    zdffqrb DNT_DW13_Q_reg_4 ( .CK(DNT_DW13_n126), .D(ADI[4]), .R(TRST_), .Q(
        DW13[4]) );
    zdffqrb DNT_DW13_Q_reg_3 ( .CK(DNT_DW13_n126), .D(ADI[3]), .R(TRST_), .Q(
        DW13[3]) );
    zdffqrb DNT_DW13_Q_reg_2 ( .CK(DNT_DW13_n126), .D(ADI[2]), .R(TRST_), .Q(
        DW13[2]) );
    zdffqrb DNT_DW13_Q_reg_1 ( .CK(DNT_DW13_n126), .D(ADI[1]), .R(TRST_), .Q(
        DW13[1]) );
    zdffqrb DNT_DW13_Q_reg_0 ( .CK(DNT_DW13_n126), .D(ADI[0]), .R(TRST_), .Q(
        DW13[0]) );
    zbfb DNT_DW13_U80 ( .A(FLOPS_CLK_13), .Y(DNT_DW13_n126) );
    zbfb DNT_DW13_U81 ( .A(FLOPS_CLK_13), .Y(DNT_DW13_n127) );
    zdffqrb DNT_DW3_Q_reg_31 ( .CK(DNT_DW3_n127), .D(AD3IN_31), .R(TRST_), .Q(
        DW3[31]) );
    zdffqrb DNT_DW3_Q_reg_30 ( .CK(DNT_DW3_n127), .D(AD3IN_30), .R(TRST_), .Q(
        DW3[30]) );
    zdffqrb DNT_DW3_Q_reg_29 ( .CK(DNT_DW3_n127), .D(AD3IN_29), .R(TRST_), .Q(
        DW3[29]) );
    zdffqrb DNT_DW3_Q_reg_28 ( .CK(DNT_DW3_n127), .D(AD3IN_28), .R(TRST_), .Q(
        DW3[28]) );
    zdffqrb DNT_DW3_Q_reg_27 ( .CK(DNT_DW3_n127), .D(AD3IN_27), .R(TRST_), .Q(
        DW3[27]) );
    zdffqrb DNT_DW3_Q_reg_26 ( .CK(DNT_DW3_n127), .D(AD3IN_26), .R(TRST_), .Q(
        DW3[26]) );
    zdffqrb DNT_DW3_Q_reg_25 ( .CK(DNT_DW3_n127), .D(AD3IN_25), .R(TRST_), .Q(
        DW3[25]) );
    zdffqrb DNT_DW3_Q_reg_24 ( .CK(DNT_DW3_n127), .D(AD3IN_24), .R(TRST_), .Q(
        DW3[24]) );
    zdffqrb DNT_DW3_Q_reg_23 ( .CK(DNT_DW3_n127), .D(AD3IN_23), .R(TRST_), .Q(
        DW3[23]) );
    zdffqrb DNT_DW3_Q_reg_22 ( .CK(DNT_DW3_n127), .D(AD3IN_22), .R(TRST_), .Q(
        DW3[22]) );
    zdffqrb DNT_DW3_Q_reg_21 ( .CK(DNT_DW3_n127), .D(AD3IN_21), .R(TRST_), .Q(
        DW3[21]) );
    zdffqrb DNT_DW3_Q_reg_20 ( .CK(DNT_DW3_n127), .D(AD3IN_20), .R(TRST_), .Q(
        DW3[20]) );
    zdffqrb DNT_DW3_Q_reg_19 ( .CK(DNT_DW3_n127), .D(AD3IN_19), .R(TRST_), .Q(
        DW3[19]) );
    zdffqrb DNT_DW3_Q_reg_18 ( .CK(DNT_DW3_n127), .D(AD3IN_18), .R(TRST_), .Q(
        DW3[18]) );
    zdffqrb DNT_DW3_Q_reg_17 ( .CK(DNT_DW3_n127), .D(AD3IN_17), .R(TRST_), .Q(
        DW3[17]) );
    zdffqrb DNT_DW3_Q_reg_16 ( .CK(DNT_DW3_n127), .D(AD3IN_16), .R(TRST_), .Q(
        DW3[16]) );
    zdffqrb DNT_DW3_Q_reg_15 ( .CK(DNT_DW3_n126), .D(AD3IN_15), .R(TRST_), .Q(
        DW3[15]) );
    zdffqrb DNT_DW3_Q_reg_14 ( .CK(DNT_DW3_n126), .D(AD3IN_14), .R(TRST_), .Q(
        DW3[14]) );
    zdffqrb DNT_DW3_Q_reg_13 ( .CK(DNT_DW3_n126), .D(AD3IN_13), .R(TRST_), .Q(
        DW3[13]) );
    zdffqrb DNT_DW3_Q_reg_12 ( .CK(DNT_DW3_n126), .D(AD3IN_12), .R(TRST_), .Q(
        DW3[12]) );
    zdffqrb DNT_DW3_Q_reg_11 ( .CK(DNT_DW3_n126), .D(AD3IN_11), .R(TRST_), .Q(
        DW3[11]) );
    zdffqrb DNT_DW3_Q_reg_10 ( .CK(DNT_DW3_n126), .D(AD3IN_10), .R(TRST_), .Q(
        DW3[10]) );
    zdffqrb DNT_DW3_Q_reg_9 ( .CK(DNT_DW3_n126), .D(AD3IN_9), .R(TRST_), .Q(
        DW3[9]) );
    zdffqrb DNT_DW3_Q_reg_8 ( .CK(DNT_DW3_n126), .D(AD3IN_8), .R(TRST_), .Q(
        DW3[8]) );
    zdffqrb DNT_DW3_Q_reg_7 ( .CK(DNT_DW3_n126), .D(AD3IN_7), .R(TRST_), .Q(
        DW3[7]) );
    zdffqrb DNT_DW3_Q_reg_6 ( .CK(DNT_DW3_n126), .D(AD3IN_6), .R(TRST_), .Q(
        DW3[6]) );
    zdffqrb DNT_DW3_Q_reg_5 ( .CK(DNT_DW3_n126), .D(AD3IN_5), .R(TRST_), .Q(
        DW3[5]) );
    zdffqrb DNT_DW3_Q_reg_4 ( .CK(DNT_DW3_n126), .D(AD3IN_4), .R(TRST_), .Q(
        DW3[4]) );
    zdffqrb DNT_DW3_Q_reg_3 ( .CK(DNT_DW3_n126), .D(AD3IN_3), .R(TRST_), .Q(
        DW3[3]) );
    zdffqrb DNT_DW3_Q_reg_2 ( .CK(DNT_DW3_n126), .D(AD3IN_2), .R(TRST_), .Q(
        DW3[2]) );
    zdffqrb DNT_DW3_Q_reg_1 ( .CK(DNT_DW3_n126), .D(AD3IN_1), .R(TRST_), .Q(
        DW3[1]) );
    zdffqrb DNT_DW3_Q_reg_0 ( .CK(DNT_DW3_n126), .D(AD3IN_0), .R(TRST_), .Q(
        DW3[0]) );
    zbfb DNT_DW3_U80 ( .A(FLOPS_CLK_3), .Y(DNT_DW3_n126) );
    zbfb DNT_DW3_U81 ( .A(FLOPS_CLK_3), .Y(DNT_DW3_n127) );
    zdffqrb DNT_DW12_Q_reg_31 ( .CK(DNT_DW12_n127), .D(ADI[31]), .R(TRST_), 
        .Q(DW12[31]) );
    zdffqrb DNT_DW12_Q_reg_30 ( .CK(DNT_DW12_n127), .D(ADI[30]), .R(TRST_), 
        .Q(DW12[30]) );
    zdffqrb DNT_DW12_Q_reg_29 ( .CK(DNT_DW12_n127), .D(ADI[29]), .R(TRST_), 
        .Q(DW12[29]) );
    zdffqrb DNT_DW12_Q_reg_28 ( .CK(DNT_DW12_n127), .D(ADI[28]), .R(TRST_), 
        .Q(DW12[28]) );
    zdffqrb DNT_DW12_Q_reg_27 ( .CK(DNT_DW12_n127), .D(ADI[27]), .R(TRST_), 
        .Q(DW12[27]) );
    zdffqrb DNT_DW12_Q_reg_26 ( .CK(DNT_DW12_n127), .D(ADI[26]), .R(TRST_), 
        .Q(DW12[26]) );
    zdffqrb DNT_DW12_Q_reg_25 ( .CK(DNT_DW12_n127), .D(ADI[25]), .R(TRST_), 
        .Q(DW12[25]) );
    zdffqrb DNT_DW12_Q_reg_24 ( .CK(DNT_DW12_n127), .D(ADI[24]), .R(TRST_), 
        .Q(DW12[24]) );
    zdffqrb DNT_DW12_Q_reg_23 ( .CK(DNT_DW12_n127), .D(ADI[23]), .R(TRST_), 
        .Q(DW12[23]) );
    zdffqrb DNT_DW12_Q_reg_22 ( .CK(DNT_DW12_n127), .D(ADI[22]), .R(TRST_), 
        .Q(DW12[22]) );
    zdffqrb DNT_DW12_Q_reg_21 ( .CK(DNT_DW12_n127), .D(ADI[21]), .R(TRST_), 
        .Q(DW12[21]) );
    zdffqrb DNT_DW12_Q_reg_20 ( .CK(DNT_DW12_n127), .D(ADI[20]), .R(TRST_), 
        .Q(DW12[20]) );
    zdffqrb DNT_DW12_Q_reg_19 ( .CK(DNT_DW12_n127), .D(ADI[19]), .R(TRST_), 
        .Q(DW12[19]) );
    zdffqrb DNT_DW12_Q_reg_18 ( .CK(DNT_DW12_n127), .D(ADI[18]), .R(TRST_), 
        .Q(DW12[18]) );
    zdffqrb DNT_DW12_Q_reg_17 ( .CK(DNT_DW12_n127), .D(ADI[17]), .R(TRST_), 
        .Q(DW12[17]) );
    zdffqrb DNT_DW12_Q_reg_16 ( .CK(DNT_DW12_n127), .D(ADI[16]), .R(TRST_), 
        .Q(DW12[16]) );
    zdffqrb DNT_DW12_Q_reg_15 ( .CK(DNT_DW12_n126), .D(ADI[15]), .R(TRST_), 
        .Q(DW12[15]) );
    zdffqrb DNT_DW12_Q_reg_14 ( .CK(DNT_DW12_n126), .D(ADI[14]), .R(TRST_), 
        .Q(DW12[14]) );
    zdffqrb DNT_DW12_Q_reg_13 ( .CK(DNT_DW12_n126), .D(ADI[13]), .R(TRST_), 
        .Q(DW12[13]) );
    zdffqrb DNT_DW12_Q_reg_12 ( .CK(DNT_DW12_n126), .D(ADI[12]), .R(TRST_), 
        .Q(DW12[12]) );
    zdffqrb DNT_DW12_Q_reg_11 ( .CK(DNT_DW12_n126), .D(ADI[11]), .R(TRST_), 
        .Q(DW12[11]) );
    zdffqrb DNT_DW12_Q_reg_10 ( .CK(DNT_DW12_n126), .D(ADI[10]), .R(TRST_), 
        .Q(DW12[10]) );
    zdffqrb DNT_DW12_Q_reg_9 ( .CK(DNT_DW12_n126), .D(ADI[9]), .R(TRST_), .Q(
        DW12[9]) );
    zdffqrb DNT_DW12_Q_reg_8 ( .CK(DNT_DW12_n126), .D(ADI[8]), .R(TRST_), .Q(
        DW12[8]) );
    zdffqrb DNT_DW12_Q_reg_7 ( .CK(DNT_DW12_n126), .D(ADI[7]), .R(TRST_), .Q(
        DW12[7]) );
    zdffqrb DNT_DW12_Q_reg_6 ( .CK(DNT_DW12_n126), .D(ADI[6]), .R(TRST_), .Q(
        DW12[6]) );
    zdffqrb DNT_DW12_Q_reg_5 ( .CK(DNT_DW12_n126), .D(ADI[5]), .R(TRST_), .Q(
        DW12[5]) );
    zdffqrb DNT_DW12_Q_reg_4 ( .CK(DNT_DW12_n126), .D(ADI[4]), .R(TRST_), .Q(
        DW12[4]) );
    zdffqrb DNT_DW12_Q_reg_3 ( .CK(DNT_DW12_n126), .D(ADI[3]), .R(TRST_), .Q(
        DW12[3]) );
    zdffqrb DNT_DW12_Q_reg_2 ( .CK(DNT_DW12_n126), .D(ADI[2]), .R(TRST_), .Q(
        DW12[2]) );
    zdffqrb DNT_DW12_Q_reg_1 ( .CK(DNT_DW12_n126), .D(ADI[1]), .R(TRST_), .Q(
        DW12[1]) );
    zdffqrb DNT_DW12_Q_reg_0 ( .CK(DNT_DW12_n126), .D(ADI[0]), .R(TRST_), .Q(
        DW12[0]) );
    zbfb DNT_DW12_U80 ( .A(FLOPS_CLK_12), .Y(DNT_DW12_n126) );
    zbfb DNT_DW12_U81 ( .A(FLOPS_CLK_12), .Y(DNT_DW12_n127) );
    zdffqrb DNT_DW4_Q_reg_31 ( .CK(DNT_DW4_n127), .D(AD4IN_31), .R(TRST_), .Q(
        DW4[31]) );
    zdffqrb DNT_DW4_Q_reg_30 ( .CK(DNT_DW4_n127), .D(AD4IN_30), .R(TRST_), .Q(
        DW4[30]) );
    zdffqrb DNT_DW4_Q_reg_29 ( .CK(DNT_DW4_n127), .D(AD4IN_29), .R(TRST_), .Q(
        DW4[29]) );
    zdffqrb DNT_DW4_Q_reg_28 ( .CK(DNT_DW4_n127), .D(AD4IN_28), .R(TRST_), .Q(
        DW4[28]) );
    zdffqrb DNT_DW4_Q_reg_27 ( .CK(DNT_DW4_n127), .D(AD4IN_27), .R(TRST_), .Q(
        DW4[27]) );
    zdffqrb DNT_DW4_Q_reg_26 ( .CK(DNT_DW4_n127), .D(AD4IN_26), .R(TRST_), .Q(
        DW4[26]) );
    zdffqrb DNT_DW4_Q_reg_25 ( .CK(DNT_DW4_n127), .D(AD4IN_25), .R(TRST_), .Q(
        DW4[25]) );
    zdffqrb DNT_DW4_Q_reg_24 ( .CK(DNT_DW4_n127), .D(AD4IN_24), .R(TRST_), .Q(
        DW4[24]) );
    zdffqrb DNT_DW4_Q_reg_23 ( .CK(DNT_DW4_n127), .D(AD4IN_23), .R(TRST_), .Q(
        DW4[23]) );
    zdffqrb DNT_DW4_Q_reg_22 ( .CK(DNT_DW4_n127), .D(AD4IN_22), .R(TRST_), .Q(
        DW4[22]) );
    zdffqrb DNT_DW4_Q_reg_21 ( .CK(DNT_DW4_n127), .D(AD4IN_21), .R(TRST_), .Q(
        DW4[21]) );
    zdffqrb DNT_DW4_Q_reg_20 ( .CK(DNT_DW4_n127), .D(AD4IN_20), .R(TRST_), .Q(
        DW4[20]) );
    zdffqrb DNT_DW4_Q_reg_19 ( .CK(DNT_DW4_n127), .D(AD4IN_19), .R(TRST_), .Q(
        DW4[19]) );
    zdffqrb DNT_DW4_Q_reg_18 ( .CK(DNT_DW4_n127), .D(AD4IN_18), .R(TRST_), .Q(
        DW4[18]) );
    zdffqrb DNT_DW4_Q_reg_17 ( .CK(DNT_DW4_n127), .D(AD4IN_17), .R(TRST_), .Q(
        DW4[17]) );
    zdffqrb DNT_DW4_Q_reg_16 ( .CK(DNT_DW4_n127), .D(AD4IN_16), .R(TRST_), .Q(
        DW4[16]) );
    zdffqrb DNT_DW4_Q_reg_15 ( .CK(DNT_DW4_n126), .D(AD4IN_15), .R(TRST_), .Q(
        DW4[15]) );
    zdffqrb DNT_DW4_Q_reg_14 ( .CK(DNT_DW4_n126), .D(AD4IN_14), .R(TRST_), .Q(
        DW4[14]) );
    zdffqrb DNT_DW4_Q_reg_13 ( .CK(DNT_DW4_n126), .D(AD4IN_13), .R(TRST_), .Q(
        DW4[13]) );
    zdffqrb DNT_DW4_Q_reg_12 ( .CK(DNT_DW4_n126), .D(AD4IN_12), .R(TRST_), .Q(
        DW4[12]) );
    zdffqrb DNT_DW4_Q_reg_11 ( .CK(DNT_DW4_n126), .D(AD4IN_11), .R(TRST_), .Q(
        DW4[11]) );
    zdffqrb DNT_DW4_Q_reg_10 ( .CK(DNT_DW4_n126), .D(AD4IN_10), .R(TRST_), .Q(
        DW4[10]) );
    zdffqrb DNT_DW4_Q_reg_9 ( .CK(DNT_DW4_n126), .D(AD4IN_9), .R(TRST_), .Q(
        DW4[9]) );
    zdffqrb DNT_DW4_Q_reg_8 ( .CK(DNT_DW4_n126), .D(AD4IN_8), .R(TRST_), .Q(
        DW4[8]) );
    zdffqrb DNT_DW4_Q_reg_7 ( .CK(DNT_DW4_n126), .D(AD4IN_7), .R(TRST_), .Q(
        DW4[7]) );
    zdffqrb DNT_DW4_Q_reg_6 ( .CK(DNT_DW4_n126), .D(AD4IN_6), .R(TRST_), .Q(
        DW4[6]) );
    zdffqrb DNT_DW4_Q_reg_5 ( .CK(DNT_DW4_n126), .D(AD4IN_5), .R(TRST_), .Q(
        DW4[5]) );
    zdffqrb DNT_DW4_Q_reg_4 ( .CK(DNT_DW4_n126), .D(AD4IN_4), .R(TRST_), .Q(
        DW4[4]) );
    zdffqrb DNT_DW4_Q_reg_3 ( .CK(DNT_DW4_n126), .D(AD4IN_3), .R(TRST_), .Q(
        DW4[3]) );
    zdffqrb DNT_DW4_Q_reg_2 ( .CK(DNT_DW4_n126), .D(AD4IN_2), .R(TRST_), .Q(
        DW4[2]) );
    zdffqrb DNT_DW4_Q_reg_1 ( .CK(DNT_DW4_n126), .D(AD4IN_1), .R(TRST_), .Q(
        DW4[1]) );
    zdffqrb DNT_DW4_Q_reg_0 ( .CK(DNT_DW4_n126), .D(AD4IN_0), .R(TRST_), .Q(
        DW4[0]) );
    zbfb DNT_DW4_U80 ( .A(FLOPS_CLK_4), .Y(DNT_DW4_n126) );
    zbfb DNT_DW4_U81 ( .A(FLOPS_CLK_4), .Y(DNT_DW4_n127) );
    zdffqrb DNT_DW15_Q_reg_31 ( .CK(DNT_DW15_n127), .D(n445), .R(TRST_), .Q(
        DW15[31]) );
    zdffqrb DNT_DW15_Q_reg_30 ( .CK(DNT_DW15_n127), .D(n470), .R(TRST_), .Q(
        DW15[30]) );
    zdffqrb DNT_DW15_Q_reg_29 ( .CK(DNT_DW15_n127), .D(n475), .R(TRST_), .Q(
        DW15[29]) );
    zdffqrb DNT_DW15_Q_reg_28 ( .CK(DNT_DW15_n127), .D(n453), .R(TRST_), .Q(
        DW15[28]) );
    zdffqrb DNT_DW15_Q_reg_27 ( .CK(DNT_DW15_n127), .D(n465), .R(TRST_), .Q(
        DW15[27]) );
    zdffqrb DNT_DW15_Q_reg_26 ( .CK(DNT_DW15_n127), .D(n459), .R(TRST_), .Q(
        DW15[26]) );
    zdffqrb DNT_DW15_Q_reg_25 ( .CK(DNT_DW15_n127), .D(n464), .R(TRST_), .Q(
        DW15[25]) );
    zdffqrb DNT_DW15_Q_reg_24 ( .CK(DNT_DW15_n127), .D(n456), .R(TRST_), .Q(
        DW15[24]) );
    zdffqrb DNT_DW15_Q_reg_23 ( .CK(DNT_DW15_n127), .D(n449), .R(TRST_), .Q(
        DW15[23]) );
    zdffqrb DNT_DW15_Q_reg_22 ( .CK(DNT_DW15_n127), .D(n468), .R(TRST_), .Q(
        DW15[22]) );
    zdffqrb DNT_DW15_Q_reg_21 ( .CK(DNT_DW15_n127), .D(n457), .R(TRST_), .Q(
        DW15[21]) );
    zdffqrb DNT_DW15_Q_reg_20 ( .CK(DNT_DW15_n127), .D(n476), .R(TRST_), .Q(
        DW15[20]) );
    zdffqrb DNT_DW15_Q_reg_19 ( .CK(DNT_DW15_n127), .D(n466), .R(TRST_), .Q(
        DW15[19]) );
    zdffqrb DNT_DW15_Q_reg_18 ( .CK(DNT_DW15_n127), .D(n452), .R(TRST_), .Q(
        DW15[18]) );
    zdffqrb DNT_DW15_Q_reg_17 ( .CK(DNT_DW15_n127), .D(n472), .R(TRST_), .Q(
        DW15[17]) );
    zdffqrb DNT_DW15_Q_reg_16 ( .CK(DNT_DW15_n127), .D(n446), .R(TRST_), .Q(
        DW15[16]) );
    zdffqrb DNT_DW15_Q_reg_15 ( .CK(DNT_DW15_n126), .D(n471), .R(TRST_), .Q(
        DW15[15]) );
    zdffqrb DNT_DW15_Q_reg_14 ( .CK(DNT_DW15_n126), .D(n455), .R(TRST_), .Q(
        DW15[14]) );
    zdffqrb DNT_DW15_Q_reg_13 ( .CK(DNT_DW15_n126), .D(n461), .R(TRST_), .Q(
        DW15[13]) );
    zdffqrb DNT_DW15_Q_reg_12 ( .CK(DNT_DW15_n126), .D(n469), .R(TRST_), .Q(
        DW15[12]) );
    zdffqrb DNT_DW15_Q_reg_11 ( .CK(DNT_DW15_n126), .D(n448), .R(TRST_), .Q(
        DW15[11]) );
    zdffqrb DNT_DW15_Q_reg_10 ( .CK(DNT_DW15_n126), .D(n460), .R(TRST_), .Q(
        DW15[10]) );
    zdffqrb DNT_DW15_Q_reg_9 ( .CK(DNT_DW15_n126), .D(n454), .R(TRST_), .Q(
        DW15[9]) );
    zdffqrb DNT_DW15_Q_reg_8 ( .CK(DNT_DW15_n126), .D(n462), .R(TRST_), .Q(
        DW15[8]) );
    zdffqrb DNT_DW15_Q_reg_7 ( .CK(DNT_DW15_n126), .D(n447), .R(TRST_), .Q(
        DW15[7]) );
    zdffqrb DNT_DW15_Q_reg_6 ( .CK(DNT_DW15_n126), .D(n474), .R(TRST_), .Q(
        DW15[6]) );
    zdffqrb DNT_DW15_Q_reg_5 ( .CK(DNT_DW15_n126), .D(n451), .R(TRST_), .Q(
        DW15[5]) );
    zdffqrb DNT_DW15_Q_reg_4 ( .CK(DNT_DW15_n126), .D(n473), .R(TRST_), .Q(
        DW15[4]) );
    zdffqrb DNT_DW15_Q_reg_3 ( .CK(DNT_DW15_n126), .D(n467), .R(TRST_), .Q(
        DW15[3]) );
    zdffqrb DNT_DW15_Q_reg_2 ( .CK(DNT_DW15_n126), .D(n463), .R(TRST_), .Q(
        DW15[2]) );
    zdffqrb DNT_DW15_Q_reg_1 ( .CK(DNT_DW15_n126), .D(n458), .R(TRST_), .Q(
        DW15[1]) );
    zdffqrb DNT_DW15_Q_reg_0 ( .CK(DNT_DW15_n126), .D(n450), .R(TRST_), .Q(
        DW15[0]) );
    zbfb DNT_DW15_U80 ( .A(FLOPS_CLK_15), .Y(DNT_DW15_n126) );
    zbfb DNT_DW15_U81 ( .A(FLOPS_CLK_15), .Y(DNT_DW15_n127) );
endmodule


module ASYNC_CACHE ( LDW, ADI, PCICLK, TRST_, CACHE_EN, DW0, DW1, DW2, DW3, 
    DW4, DW5, DW6, DW7, DW8, DW9, DW10, DW11, CACHEPHASE, UP_DW3, UP_DW5, 
    UP_DW6, UP_DW7, UP_LDW3, UP_LDW5, UP_LDW6, UP_LDW7, ATPG_ENI );
input  [15:0] LDW;
output [31:0] DW0;
input  [31:0] ADI;
output [31:0] DW7;
output [31:0] DW9;
input  [31:0] UP_DW6;
output [31:0] DW1;
output [31:0] DW6;
input  [31:0] UP_DW7;
output [31:0] DW2;
output [31:0] DW3;
output [31:0] DW8;
output [31:0] DW4;
input  [31:0] UP_DW5;
output [31:0] DW5;
output [31:0] DW10;
output [31:0] DW11;
input  [31:0] UP_DW3;
input  PCICLK, TRST_, CACHE_EN, CACHEPHASE, UP_LDW3, UP_LDW5, UP_LDW6, UP_LDW7, 
    ATPG_ENI;
    wire AD5IN_3, FLOPS_CLK_11, AD6IN_9, AD3IN_25, n_16, AD3IN_2, AD7IN_21, 
        AD7IN_5, AD6IN_13, AD5IN_10, AD3IN_19, n_23, AD6IN_0, AD5IN_25, 
        AD7IN_28, AD6IN_26, AD7IN_14, AD5IN_19, n_18, AD3IN_10, AD3IN_30, 
        AD3IN_17, AD7IN_13, AD6IN_21, AD5IN_22, n_9, n_11, n_24, AD6IN_7, 
        FLOPS_CLK_13, AD6IN_28, AD5IN_30, AD5IN_17, AD3IN_5, AD6IN_14, AD7IN_2, 
        AD7IN_26, AD5IN_4, AD3IN_22, FLOPS_CLK_4, AD6IN_6, FLOPS_CLK_12, 
        AD5IN_23, n_19, AD7IN_12, AD6IN_20, AD3IN_31, AD3IN_16, AD5IN_5, n_10, 
        AD3IN_23, FLOPS_CLK_5, AD3IN_4, AD6IN_15, AD7IN_3, AD7IN_27, AD6IN_29, 
        AD5IN_31, AD5IN_16, AD3IN_18, AD5IN_11, AD3IN_3, AD7IN_20, AD7IN_4, 
        AD6IN_12, AD5IN_2, AD6IN_8, AD3IN_24, FLOPS_CLK_10, AD3IN_11, AD6IN_27, 
        AD7IN_15, n_22, AD5IN_18, AD5IN_24, AD7IN_29, AD6IN_1, FLOPS_CLK_8, 
        AD3IN_26, AD5IN_0, FLOPS_CLK_14, AD7IN_6, AD7IN_22, AD6IN_10, AD3IN_1, 
        AD5IN_13, n_20, AD6IN_3, AD5IN_9, AD6IN_19, AD3IN_8, AD5IN_26, 
        AD7IN_17, AD6IN_25, AD7IN_30, AD3IN_13, AD3IN_14, AD6IN_22, AD7IN_10, 
        AD7IN_8, n_12, AD5IN_21, AD3IN_28, AD6IN_4, AD5IN_14, AD7IN_19, 
        AD6IN_30, AD7IN_25, AD6IN_17, AD7IN_1, AD5IN_28, AD3IN_21, AD3IN_6, 
        FLOPS_CLK_7, AD5IN_7, AD3IN_29, AD6IN_5, AD7IN_9, AD5IN_20, AD6IN_23, 
        AD7IN_11, AD3IN_20, AD3IN_15, FLOPS_CLK_6, AD5IN_6, AD6IN_31, AD7IN_24, 
        AD6IN_16, AD7IN_0, AD5IN_29, AD3IN_7, AD5IN_15, AD7IN_18, AD5IN_12, 
        AD7IN_7, AD6IN_11, AD7IN_23, AD3IN_0, AD3IN_27, FLOPS_CLK_9, AD5IN_1, 
        FLOPS_CLK_15, AD3IN_12, n_21, AD7IN_16, AD6IN_24, AD7IN_31, AD6IN_18, 
        AD3IN_9, AD5IN_27, AD6IN_2, AD5IN_8, n267, n268, n269, n270, n271, 
        n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
        n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
        n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
        n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
        n320, n321, n322, DNT_DW6_n126, DNT_DW6_n127, DNT_DW1_n126, 
        DNT_DW1_n127, DNT_DW10_n126, DNT_DW10_n127, DNT_DW8_n126, DNT_DW8_n127, 
        DNT_DW0_n126, DNT_DW0_n127, DNT_DW11_n126, DNT_DW11_n127, DNT_DW9_n126, 
        DNT_DW9_n127, DNT_DW7_n126, DNT_DW7_n127, DNT_DW5_n126, DNT_DW5_n127, 
        DNT_DW2_n126, DNT_DW2_n127, DNT_DW3_n126, DNT_DW3_n127, DNT_DW4_n126, 
        DNT_DW4_n127;
    zan2b U40 ( .A(LDW[4]), .B(n321), .Y(n_16) );
    zan2b U41 ( .A(LDW[2]), .B(n321), .Y(n_18) );
    zan2b U42 ( .A(CACHE_EN), .B(LDW[11]), .Y(n_9) );
    zan2b U43 ( .A(LDW[0]), .B(n321), .Y(n_20) );
    zan2b U44 ( .A(LDW[8]), .B(n321), .Y(n_12) );
    zan2b U45 ( .A(LDW[10]), .B(n321), .Y(n_10) );
    zao21b U46 ( .A(UP_DW3[0]), .B(n304), .C(n298), .Y(AD3IN_0) );
    zao21b U47 ( .A(UP_DW3[1]), .B(n312), .C(n297), .Y(AD3IN_1) );
    zao21b U48 ( .A(UP_DW3[3]), .B(n314), .C(n295), .Y(AD3IN_3) );
    zao21b U49 ( .A(UP_DW3[4]), .B(n304), .C(n294), .Y(AD3IN_4) );
    zao21b U50 ( .A(UP_DW3[5]), .B(n305), .C(n293), .Y(AD3IN_5) );
    zao21b U51 ( .A(UP_DW3[6]), .B(n310), .C(n292), .Y(AD3IN_6) );
    zao21b U52 ( .A(UP_DW3[7]), .B(n314), .C(n291), .Y(AD3IN_7) );
    zao21b U53 ( .A(UP_DW3[9]), .B(n313), .C(n289), .Y(AD3IN_9) );
    zao21b U54 ( .A(UP_DW3[11]), .B(n304), .C(n287), .Y(AD3IN_11) );
    zao21b U55 ( .A(UP_DW3[12]), .B(n305), .C(n286), .Y(AD3IN_12) );
    zao21b U56 ( .A(UP_DW3[13]), .B(n312), .C(n285), .Y(AD3IN_13) );
    zao21b U57 ( .A(UP_DW3[15]), .B(n314), .C(n283), .Y(AD3IN_15) );
    zao21b U58 ( .A(UP_DW3[18]), .B(n309), .C(n280), .Y(AD3IN_18) );
    zao21b U59 ( .A(UP_DW3[19]), .B(n305), .C(n279), .Y(AD3IN_19) );
    zao21b U60 ( .A(UP_DW3[22]), .B(n313), .C(n276), .Y(AD3IN_22) );
    zao21b U61 ( .A(UP_DW3[23]), .B(n312), .C(n275), .Y(AD3IN_23) );
    zao21b U62 ( .A(UP_DW3[24]), .B(n299), .C(n274), .Y(AD3IN_24) );
    zao21b U63 ( .A(UP_DW3[28]), .B(n313), .C(n270), .Y(AD3IN_28) );
    zao21b U64 ( .A(UP_DW3[30]), .B(n314), .C(n268), .Y(AD3IN_30) );
    zao21b U65 ( .A(UP_DW3[31]), .B(n302), .C(n267), .Y(AD3IN_31) );
    zao21b U66 ( .A(UP_DW5[1]), .B(n302), .C(n297), .Y(AD5IN_1) );
    zao21b U67 ( .A(UP_DW5[2]), .B(n307), .C(n296), .Y(AD5IN_2) );
    zao21b U68 ( .A(UP_DW5[4]), .B(n302), .C(n294), .Y(AD5IN_4) );
    zao21b U69 ( .A(UP_DW5[6]), .B(n301), .C(n292), .Y(AD5IN_6) );
    zao21b U70 ( .A(UP_DW5[7]), .B(n308), .C(n291), .Y(AD5IN_7) );
    zao21b U71 ( .A(UP_DW5[10]), .B(n307), .C(n288), .Y(AD5IN_10) );
    zao21b U72 ( .A(UP_DW5[15]), .B(n317), .C(n283), .Y(AD5IN_15) );
    zao21b U73 ( .A(UP_DW5[18]), .B(n318), .C(n280), .Y(AD5IN_18) );
    zao21b U74 ( .A(UP_DW5[21]), .B(n316), .C(n277), .Y(AD5IN_21) );
    zao21b U75 ( .A(UP_DW5[23]), .B(n308), .C(n275), .Y(AD5IN_23) );
    zao21b U76 ( .A(UP_DW5[24]), .B(n319), .C(n274), .Y(AD5IN_24) );
    zao21b U77 ( .A(UP_DW5[25]), .B(n318), .C(n273), .Y(AD5IN_25) );
    zao21b U78 ( .A(UP_DW5[26]), .B(n302), .C(n272), .Y(AD5IN_26) );
    zao21b U79 ( .A(UP_DW5[29]), .B(n307), .C(n269), .Y(AD5IN_29) );
    zao21b U80 ( .A(UP_DW5[30]), .B(n317), .C(n268), .Y(AD5IN_30) );
    zao21b U81 ( .A(UP_DW7[1]), .B(n307), .C(n297), .Y(AD7IN_1) );
    zao21b U82 ( .A(UP_DW7[2]), .B(n319), .C(n296), .Y(AD7IN_2) );
    zao21b U83 ( .A(UP_DW7[5]), .B(n309), .C(n293), .Y(AD7IN_5) );
    zao21b U84 ( .A(UP_DW7[10]), .B(n318), .C(n288), .Y(AD7IN_10) );
    zao21b U85 ( .A(UP_DW7[12]), .B(n302), .C(n286), .Y(AD7IN_12) );
    zao21b U86 ( .A(UP_DW7[13]), .B(n318), .C(n285), .Y(AD7IN_13) );
    zao21b U87 ( .A(UP_DW7[14]), .B(n308), .C(n284), .Y(AD7IN_14) );
    zao21b U88 ( .A(UP_DW7[15]), .B(n308), .C(n283), .Y(AD7IN_15) );
    zao21b U89 ( .A(UP_DW7[17]), .B(n301), .C(n281), .Y(AD7IN_17) );
    zao21b U90 ( .A(UP_DW7[18]), .B(n304), .C(n280), .Y(AD7IN_18) );
    zao21b U91 ( .A(UP_DW7[22]), .B(n308), .C(n276), .Y(AD7IN_22) );
    zao21b U92 ( .A(UP_DW7[23]), .B(n316), .C(n275), .Y(AD7IN_23) );
    zao21b U93 ( .A(UP_DW7[24]), .B(n319), .C(n274), .Y(AD7IN_24) );
    zao21b U94 ( .A(UP_DW7[25]), .B(n301), .C(n273), .Y(AD7IN_25) );
    zao21b U95 ( .A(UP_DW7[26]), .B(n301), .C(n272), .Y(AD7IN_26) );
    zao21b U96 ( .A(UP_DW7[28]), .B(n316), .C(n270), .Y(AD7IN_28) );
    zao21b U97 ( .A(UP_DW7[29]), .B(n318), .C(n269), .Y(AD7IN_29) );
    zao21b U98 ( .A(UP_DW7[30]), .B(n316), .C(n268), .Y(AD7IN_30) );
    zao21b U99 ( .A(UP_DW6[1]), .B(n319), .C(n297), .Y(AD6IN_1) );
    zao21b U100 ( .A(UP_DW6[2]), .B(n314), .C(n296), .Y(AD6IN_2) );
    zao21b U101 ( .A(UP_DW6[5]), .B(n319), .C(n293), .Y(AD6IN_5) );
    zao21b U102 ( .A(UP_DW6[7]), .B(n317), .C(n291), .Y(AD6IN_7) );
    zao21b U103 ( .A(UP_DW6[8]), .B(n299), .C(n290), .Y(AD6IN_8) );
    zao21b U104 ( .A(UP_DW6[9]), .B(n317), .C(n289), .Y(AD6IN_9) );
    zao21b U105 ( .A(UP_DW6[11]), .B(n316), .C(n287), .Y(AD6IN_11) );
    zao21b U106 ( .A(UP_DW6[13]), .B(n317), .C(n285), .Y(AD6IN_13) );
    zao21b U107 ( .A(UP_DW6[16]), .B(n313), .C(n282), .Y(AD6IN_16) );
    zao21b U108 ( .A(UP_DW6[17]), .B(n301), .C(n281), .Y(AD6IN_17) );
    zao21b U109 ( .A(UP_DW6[19]), .B(n307), .C(n279), .Y(AD6IN_19) );
    zao21b U110 ( .A(UP_DW6[22]), .B(n310), .C(n276), .Y(AD6IN_22) );
    zao21b U111 ( .A(UP_DW6[24]), .B(n309), .C(n274), .Y(AD6IN_24) );
    zao21b U112 ( .A(UP_DW6[25]), .B(n310), .C(n273), .Y(AD6IN_25) );
    zao21b U113 ( .A(UP_DW6[26]), .B(n310), .C(n272), .Y(AD6IN_26) );
    zao21b U114 ( .A(UP_DW6[27]), .B(n305), .C(n271), .Y(AD6IN_27) );
    zao21b U115 ( .A(UP_DW6[28]), .B(n312), .C(n270), .Y(AD6IN_28) );
    zao21b U116 ( .A(UP_DW6[29]), .B(n314), .C(n269), .Y(AD6IN_29) );
    zao21b U117 ( .A(UP_DW6[31]), .B(n314), .C(n267), .Y(AD6IN_31) );
    zan2b U118 ( .A(ADI[31]), .B(n306), .Y(n267) );
    zan2b U119 ( .A(ADI[30]), .B(n303), .Y(n268) );
    zan2b U120 ( .A(ADI[29]), .B(n306), .Y(n269) );
    zan2b U121 ( .A(ADI[28]), .B(n300), .Y(n270) );
    zan2b U122 ( .A(ADI[27]), .B(n320), .Y(n271) );
    zan2b U123 ( .A(ADI[26]), .B(n306), .Y(n272) );
    zan2b U124 ( .A(ADI[25]), .B(n300), .Y(n273) );
    zan2b U125 ( .A(ADI[24]), .B(n320), .Y(n274) );
    zan2b U126 ( .A(ADI[23]), .B(n320), .Y(n275) );
    zan2b U127 ( .A(ADI[22]), .B(n303), .Y(n276) );
    zan2b U128 ( .A(ADI[21]), .B(n306), .Y(n277) );
    zan2b U129 ( .A(ADI[20]), .B(n320), .Y(n278) );
    zan2b U130 ( .A(ADI[19]), .B(n300), .Y(n279) );
    zan2b U131 ( .A(ADI[18]), .B(n300), .Y(n280) );
    zan2b U132 ( .A(ADI[17]), .B(n300), .Y(n281) );
    zan2b U133 ( .A(ADI[16]), .B(n300), .Y(n282) );
    zan2b U134 ( .A(ADI[15]), .B(n320), .Y(n283) );
    zan2b U135 ( .A(ADI[14]), .B(n300), .Y(n284) );
    zan2b U136 ( .A(ADI[13]), .B(n306), .Y(n285) );
    zan2b U137 ( .A(ADI[12]), .B(n303), .Y(n286) );
    zan2b U138 ( .A(ADI[11]), .B(n306), .Y(n287) );
    zan2b U139 ( .A(ADI[10]), .B(n303), .Y(n288) );
    zan2b U140 ( .A(ADI[9]), .B(n320), .Y(n289) );
    zan2b U141 ( .A(ADI[8]), .B(n306), .Y(n290) );
    zan2b U142 ( .A(ADI[7]), .B(n306), .Y(n291) );
    zan2b U143 ( .A(ADI[6]), .B(n300), .Y(n292) );
    zan2b U144 ( .A(ADI[5]), .B(n300), .Y(n293) );
    zan2b U145 ( .A(ADI[4]), .B(n303), .Y(n294) );
    zan2b U146 ( .A(ADI[3]), .B(n306), .Y(n295) );
    zan2b U147 ( .A(ADI[2]), .B(n303), .Y(n296) );
    zan2b U148 ( .A(ADI[1]), .B(n320), .Y(n297) );
    zan2b U149 ( .A(ADI[0]), .B(n303), .Y(n298) );
    ziv11b U150 ( .A(n311), .Y(n299), .Z(n300) );
    zivb U151 ( .A(n315), .Y(n302) );
    zivb U152 ( .A(n315), .Y(n301) );
    zao21b U153 ( .A(UP_DW7[11]), .B(n316), .C(n287), .Y(AD7IN_11) );
    zao21b U154 ( .A(UP_DW5[28]), .B(n318), .C(n270), .Y(AD5IN_28) );
    zao21b U155 ( .A(UP_DW5[0]), .B(n319), .C(n298), .Y(AD5IN_0) );
    zao21b U156 ( .A(UP_DW7[19]), .B(n301), .C(n279), .Y(AD7IN_19) );
    zao21b U157 ( .A(UP_DW6[15]), .B(n308), .C(n283), .Y(AD6IN_15) );
    zao21b U158 ( .A(UP_DW6[3]), .B(n302), .C(n295), .Y(AD6IN_3) );
    zao21b U159 ( .A(UP_DW5[27]), .B(n307), .C(n271), .Y(AD5IN_27) );
    zao21b U160 ( .A(UP_DW7[31]), .B(n317), .C(n267), .Y(AD7IN_31) );
    zao21b U161 ( .A(LDW[5]), .B(n321), .C(UP_LDW5), .Y(n_23) );
    zao21b U162 ( .A(LDW[7]), .B(n321), .C(UP_LDW7), .Y(n_21) );
    zao21b U163 ( .A(LDW[3]), .B(n321), .C(UP_LDW3), .Y(n_24) );
    zao21b U164 ( .A(LDW[6]), .B(n321), .C(UP_LDW6), .Y(n_22) );
    zan2b U165 ( .A(LDW[9]), .B(CACHE_EN), .Y(n_11) );
    zan2b U166 ( .A(LDW[1]), .B(CACHE_EN), .Y(n_19) );
    zivb U167 ( .A(n322), .Y(n321) );
    zivb U168 ( .A(CACHE_EN), .Y(n322) );
    zivb U169 ( .A(n314), .Y(n303) );
    zivb U170 ( .A(n314), .Y(n320) );
    zivb U171 ( .A(n311), .Y(n314) );
    zivb U172 ( .A(n311), .Y(n305) );
    zivb U173 ( .A(n311), .Y(n304) );
    zao21b U174 ( .A(UP_DW7[16]), .B(n312), .C(n282), .Y(AD7IN_16) );
    zao21b U175 ( .A(UP_DW3[26]), .B(n313), .C(n272), .Y(AD3IN_26) );
    zao21b U176 ( .A(UP_DW7[8]), .B(n309), .C(n290), .Y(AD7IN_8) );
    zao21b U177 ( .A(UP_DW6[4]), .B(n304), .C(n294), .Y(AD6IN_4) );
    zao21b U178 ( .A(UP_DW6[23]), .B(n310), .C(n275), .Y(AD6IN_23) );
    zao21b U179 ( .A(UP_DW3[21]), .B(n313), .C(n277), .Y(AD3IN_21) );
    zao21b U180 ( .A(UP_DW3[17]), .B(n305), .C(n281), .Y(AD3IN_17) );
    zivb U181 ( .A(n299), .Y(n306) );
    zivb U182 ( .A(n315), .Y(n308) );
    zivb U183 ( .A(n315), .Y(n307) );
    zao21b U184 ( .A(UP_DW7[27]), .B(n307), .C(n271), .Y(AD7IN_27) );
    zao21b U185 ( .A(UP_DW5[17]), .B(n319), .C(n281), .Y(AD5IN_17) );
    zao21b U186 ( .A(UP_DW5[19]), .B(n319), .C(n279), .Y(AD5IN_19) );
    zao21b U187 ( .A(UP_DW5[3]), .B(n307), .C(n295), .Y(AD5IN_3) );
    zao21b U188 ( .A(UP_DW5[9]), .B(n301), .C(n289), .Y(AD5IN_9) );
    zao21b U189 ( .A(UP_DW7[21]), .B(n317), .C(n277), .Y(AD7IN_21) );
    zao21b U190 ( .A(UP_DW5[11]), .B(n308), .C(n287), .Y(AD5IN_11) );
    zao21b U191 ( .A(UP_DW5[5]), .B(n316), .C(n293), .Y(AD5IN_5) );
    zao21b U192 ( .A(UP_DW5[13]), .B(n301), .C(n285), .Y(AD5IN_13) );
    zao21b U193 ( .A(UP_DW5[8]), .B(n316), .C(n290), .Y(AD5IN_8) );
    zao21b U194 ( .A(UP_DW5[14]), .B(n308), .C(n284), .Y(AD5IN_14) );
    zao21b U195 ( .A(UP_DW5[16]), .B(n302), .C(n282), .Y(AD5IN_16) );
    zao21b U196 ( .A(UP_DW7[0]), .B(n318), .C(n298), .Y(AD7IN_0) );
    zao21b U197 ( .A(UP_DW5[20]), .B(n307), .C(n278), .Y(AD5IN_20) );
    zao21b U198 ( .A(UP_DW7[20]), .B(n302), .C(n278), .Y(AD7IN_20) );
    zao21b U199 ( .A(UP_DW5[22]), .B(n318), .C(n276), .Y(AD5IN_22) );
    zao21b U200 ( .A(UP_DW5[12]), .B(n317), .C(n286), .Y(AD5IN_12) );
    zivb U201 ( .A(n311), .Y(n310) );
    zivb U202 ( .A(n311), .Y(n309) );
    zao21b U203 ( .A(n304), .B(UP_DW7[9]), .C(n289), .Y(AD7IN_9) );
    zao21b U204 ( .A(UP_DW3[2]), .B(n309), .C(n296), .Y(AD3IN_2) );
    zao21b U205 ( .A(UP_DW3[25]), .B(n309), .C(n273), .Y(AD3IN_25) );
    zao21b U206 ( .A(UP_DW7[7]), .B(n310), .C(n291), .Y(AD7IN_7) );
    zao21b U207 ( .A(UP_DW3[20]), .B(n313), .C(n278), .Y(AD3IN_20) );
    zao21b U208 ( .A(UP_DW6[18]), .B(n310), .C(n280), .Y(AD6IN_18) );
    zao21b U209 ( .A(UP_DW7[4]), .B(n305), .C(n294), .Y(AD7IN_4) );
    zao21b U210 ( .A(UP_DW3[16]), .B(n313), .C(n282), .Y(AD3IN_16) );
    zao21b U211 ( .A(UP_DW3[10]), .B(n310), .C(n288), .Y(AD3IN_10) );
    zao21b U212 ( .A(UP_DW3[29]), .B(n304), .C(n269), .Y(AD3IN_29) );
    zao21b U213 ( .A(UP_DW6[21]), .B(n309), .C(n277), .Y(AD6IN_21) );
    zao21b U214 ( .A(UP_DW3[8]), .B(n312), .C(n290), .Y(AD3IN_8) );
    zao21b U215 ( .A(UP_DW7[3]), .B(n309), .C(n295), .Y(AD7IN_3) );
    zao21b U216 ( .A(UP_DW6[10]), .B(n304), .C(n288), .Y(AD6IN_10) );
    zao21b U217 ( .A(UP_DW3[27]), .B(n305), .C(n271), .Y(AD3IN_27) );
    zao21b U218 ( .A(UP_DW6[30]), .B(n305), .C(n268), .Y(AD6IN_30) );
    zao21b U219 ( .A(UP_DW6[0]), .B(n312), .C(n298), .Y(AD6IN_0) );
    zao21b U220 ( .A(UP_DW6[12]), .B(n312), .C(n286), .Y(AD6IN_12) );
    zao21b U221 ( .A(UP_DW7[6]), .B(n312), .C(n292), .Y(AD7IN_6) );
    zao21b U222 ( .A(UP_DW6[14]), .B(n309), .C(n284), .Y(AD6IN_14) );
    zao21b U223 ( .A(UP_DW6[6]), .B(n305), .C(n292), .Y(AD6IN_6) );
    zao21b U224 ( .A(UP_DW5[31]), .B(n313), .C(n267), .Y(AD5IN_31) );
    zao21b U225 ( .A(UP_DW3[14]), .B(n304), .C(n284), .Y(AD3IN_14) );
    zao21b U226 ( .A(UP_DW6[20]), .B(n310), .C(n278), .Y(AD6IN_20) );
    zivb U227 ( .A(CACHEPHASE), .Y(n311) );
    zivb U228 ( .A(n311), .Y(n312) );
    zivb U229 ( .A(n311), .Y(n313) );
    zivb U230 ( .A(CACHEPHASE), .Y(n315) );
    zivb U231 ( .A(n315), .Y(n316) );
    zivb U232 ( .A(n315), .Y(n319) );
    zivb U233 ( .A(n315), .Y(n317) );
    zivb U234 ( .A(n315), .Y(n318) );
    zmux21hd U235 ( .A(n_9), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_15) );
    zmux21hd U236 ( .A(n_10), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_14) );
    zmux21hd U237 ( .A(n_11), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_13) );
    zmux21hd U238 ( .A(n_12), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_12) );
    zmux21hd U239 ( .A(n_21), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_11) );
    zmux21hd U240 ( .A(n_22), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_10) );
    zmux21hd U241 ( .A(n_23), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_9) );
    zmux21hd U242 ( .A(n_16), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_8) );
    zmux21hd U243 ( .A(n_24), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_7) );
    zmux21hd U244 ( .A(n_18), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_6) );
    zmux21hd U245 ( .A(n_19), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_5) );
    zmux21hd U246 ( .A(n_20), .B(PCICLK), .S(ATPG_ENI), .Y(FLOPS_CLK_4) );
    zdffqrb DNT_DW6_Q_reg_31 ( .CK(DNT_DW6_n127), .D(AD6IN_31), .R(TRST_), .Q(
        DW6[31]) );
    zdffqrb DNT_DW6_Q_reg_30 ( .CK(DNT_DW6_n127), .D(AD6IN_30), .R(TRST_), .Q(
        DW6[30]) );
    zdffqrb DNT_DW6_Q_reg_29 ( .CK(DNT_DW6_n127), .D(AD6IN_29), .R(TRST_), .Q(
        DW6[29]) );
    zdffqrb DNT_DW6_Q_reg_28 ( .CK(DNT_DW6_n127), .D(AD6IN_28), .R(TRST_), .Q(
        DW6[28]) );
    zdffqrb DNT_DW6_Q_reg_27 ( .CK(DNT_DW6_n127), .D(AD6IN_27), .R(TRST_), .Q(
        DW6[27]) );
    zdffqrb DNT_DW6_Q_reg_26 ( .CK(DNT_DW6_n127), .D(AD6IN_26), .R(TRST_), .Q(
        DW6[26]) );
    zdffqrb DNT_DW6_Q_reg_25 ( .CK(DNT_DW6_n127), .D(AD6IN_25), .R(TRST_), .Q(
        DW6[25]) );
    zdffqrb DNT_DW6_Q_reg_24 ( .CK(DNT_DW6_n127), .D(AD6IN_24), .R(TRST_), .Q(
        DW6[24]) );
    zdffqrb DNT_DW6_Q_reg_23 ( .CK(DNT_DW6_n127), .D(AD6IN_23), .R(TRST_), .Q(
        DW6[23]) );
    zdffqrb DNT_DW6_Q_reg_22 ( .CK(DNT_DW6_n127), .D(AD6IN_22), .R(TRST_), .Q(
        DW6[22]) );
    zdffqrb DNT_DW6_Q_reg_21 ( .CK(DNT_DW6_n127), .D(AD6IN_21), .R(TRST_), .Q(
        DW6[21]) );
    zdffqrb DNT_DW6_Q_reg_20 ( .CK(DNT_DW6_n127), .D(AD6IN_20), .R(TRST_), .Q(
        DW6[20]) );
    zdffqrb DNT_DW6_Q_reg_19 ( .CK(DNT_DW6_n127), .D(AD6IN_19), .R(TRST_), .Q(
        DW6[19]) );
    zdffqrb DNT_DW6_Q_reg_18 ( .CK(DNT_DW6_n127), .D(AD6IN_18), .R(TRST_), .Q(
        DW6[18]) );
    zdffqrb DNT_DW6_Q_reg_17 ( .CK(DNT_DW6_n127), .D(AD6IN_17), .R(TRST_), .Q(
        DW6[17]) );
    zdffqrb DNT_DW6_Q_reg_16 ( .CK(DNT_DW6_n127), .D(AD6IN_16), .R(TRST_), .Q(
        DW6[16]) );
    zdffqrb DNT_DW6_Q_reg_15 ( .CK(DNT_DW6_n126), .D(AD6IN_15), .R(TRST_), .Q(
        DW6[15]) );
    zdffqrb DNT_DW6_Q_reg_14 ( .CK(DNT_DW6_n126), .D(AD6IN_14), .R(TRST_), .Q(
        DW6[14]) );
    zdffqrb DNT_DW6_Q_reg_13 ( .CK(DNT_DW6_n126), .D(AD6IN_13), .R(TRST_), .Q(
        DW6[13]) );
    zdffqrb DNT_DW6_Q_reg_12 ( .CK(DNT_DW6_n126), .D(AD6IN_12), .R(TRST_), .Q(
        DW6[12]) );
    zdffqrb DNT_DW6_Q_reg_11 ( .CK(DNT_DW6_n126), .D(AD6IN_11), .R(TRST_), .Q(
        DW6[11]) );
    zdffqrb DNT_DW6_Q_reg_10 ( .CK(DNT_DW6_n126), .D(AD6IN_10), .R(TRST_), .Q(
        DW6[10]) );
    zdffqrb DNT_DW6_Q_reg_9 ( .CK(DNT_DW6_n126), .D(AD6IN_9), .R(TRST_), .Q(
        DW6[9]) );
    zdffqrb DNT_DW6_Q_reg_8 ( .CK(DNT_DW6_n126), .D(AD6IN_8), .R(TRST_), .Q(
        DW6[8]) );
    zdffqrb DNT_DW6_Q_reg_7 ( .CK(DNT_DW6_n126), .D(AD6IN_7), .R(TRST_), .Q(
        DW6[7]) );
    zdffqrb DNT_DW6_Q_reg_6 ( .CK(DNT_DW6_n126), .D(AD6IN_6), .R(TRST_), .Q(
        DW6[6]) );
    zdffqrb DNT_DW6_Q_reg_5 ( .CK(DNT_DW6_n126), .D(AD6IN_5), .R(TRST_), .Q(
        DW6[5]) );
    zdffqrb DNT_DW6_Q_reg_4 ( .CK(DNT_DW6_n126), .D(AD6IN_4), .R(TRST_), .Q(
        DW6[4]) );
    zdffqrb DNT_DW6_Q_reg_3 ( .CK(DNT_DW6_n126), .D(AD6IN_3), .R(TRST_), .Q(
        DW6[3]) );
    zdffqrb DNT_DW6_Q_reg_2 ( .CK(DNT_DW6_n126), .D(AD6IN_2), .R(TRST_), .Q(
        DW6[2]) );
    zdffqrb DNT_DW6_Q_reg_1 ( .CK(DNT_DW6_n126), .D(AD6IN_1), .R(TRST_), .Q(
        DW6[1]) );
    zdffqrb DNT_DW6_Q_reg_0 ( .CK(DNT_DW6_n126), .D(AD6IN_0), .R(TRST_), .Q(
        DW6[0]) );
    zbfb DNT_DW6_U80 ( .A(FLOPS_CLK_10), .Y(DNT_DW6_n126) );
    zbfb DNT_DW6_U81 ( .A(FLOPS_CLK_10), .Y(DNT_DW6_n127) );
    zdffqrb DNT_DW1_Q_reg_31 ( .CK(DNT_DW1_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW1[31]) );
    zdffqrb DNT_DW1_Q_reg_30 ( .CK(DNT_DW1_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW1[30]) );
    zdffqrb DNT_DW1_Q_reg_29 ( .CK(DNT_DW1_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW1[29]) );
    zdffqrb DNT_DW1_Q_reg_28 ( .CK(DNT_DW1_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW1[28]) );
    zdffqrb DNT_DW1_Q_reg_27 ( .CK(DNT_DW1_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW1[27]) );
    zdffqrb DNT_DW1_Q_reg_26 ( .CK(DNT_DW1_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW1[26]) );
    zdffqrb DNT_DW1_Q_reg_25 ( .CK(DNT_DW1_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW1[25]) );
    zdffqrb DNT_DW1_Q_reg_24 ( .CK(DNT_DW1_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW1[24]) );
    zdffqrb DNT_DW1_Q_reg_23 ( .CK(DNT_DW1_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW1[23]) );
    zdffqrb DNT_DW1_Q_reg_22 ( .CK(DNT_DW1_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW1[22]) );
    zdffqrb DNT_DW1_Q_reg_21 ( .CK(DNT_DW1_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW1[21]) );
    zdffqrb DNT_DW1_Q_reg_20 ( .CK(DNT_DW1_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW1[20]) );
    zdffqrb DNT_DW1_Q_reg_19 ( .CK(DNT_DW1_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW1[19]) );
    zdffqrb DNT_DW1_Q_reg_18 ( .CK(DNT_DW1_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW1[18]) );
    zdffqrb DNT_DW1_Q_reg_17 ( .CK(DNT_DW1_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW1[17]) );
    zdffqrb DNT_DW1_Q_reg_16 ( .CK(DNT_DW1_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW1[16]) );
    zdffqrb DNT_DW1_Q_reg_15 ( .CK(DNT_DW1_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW1[15]) );
    zdffqrb DNT_DW1_Q_reg_14 ( .CK(DNT_DW1_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW1[14]) );
    zdffqrb DNT_DW1_Q_reg_13 ( .CK(DNT_DW1_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW1[13]) );
    zdffqrb DNT_DW1_Q_reg_12 ( .CK(DNT_DW1_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW1[12]) );
    zdffqrb DNT_DW1_Q_reg_11 ( .CK(DNT_DW1_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW1[11]) );
    zdffqrb DNT_DW1_Q_reg_10 ( .CK(DNT_DW1_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW1[10]) );
    zdffqrb DNT_DW1_Q_reg_9 ( .CK(DNT_DW1_n126), .D(ADI[9]), .R(TRST_), .Q(DW1
        [9]) );
    zdffqrb DNT_DW1_Q_reg_8 ( .CK(DNT_DW1_n126), .D(ADI[8]), .R(TRST_), .Q(DW1
        [8]) );
    zdffqrb DNT_DW1_Q_reg_7 ( .CK(DNT_DW1_n126), .D(ADI[7]), .R(TRST_), .Q(DW1
        [7]) );
    zdffqrb DNT_DW1_Q_reg_6 ( .CK(DNT_DW1_n126), .D(ADI[6]), .R(TRST_), .Q(DW1
        [6]) );
    zdffqrb DNT_DW1_Q_reg_5 ( .CK(DNT_DW1_n126), .D(ADI[5]), .R(TRST_), .Q(DW1
        [5]) );
    zdffqrb DNT_DW1_Q_reg_4 ( .CK(DNT_DW1_n126), .D(ADI[4]), .R(TRST_), .Q(DW1
        [4]) );
    zdffqrb DNT_DW1_Q_reg_3 ( .CK(DNT_DW1_n126), .D(ADI[3]), .R(TRST_), .Q(DW1
        [3]) );
    zdffqrb DNT_DW1_Q_reg_2 ( .CK(DNT_DW1_n126), .D(ADI[2]), .R(TRST_), .Q(DW1
        [2]) );
    zdffqrb DNT_DW1_Q_reg_1 ( .CK(DNT_DW1_n126), .D(ADI[1]), .R(TRST_), .Q(DW1
        [1]) );
    zdffqrb DNT_DW1_Q_reg_0 ( .CK(DNT_DW1_n126), .D(ADI[0]), .R(TRST_), .Q(DW1
        [0]) );
    zbfb DNT_DW1_U80 ( .A(FLOPS_CLK_5), .Y(DNT_DW1_n126) );
    zbfb DNT_DW1_U81 ( .A(FLOPS_CLK_5), .Y(DNT_DW1_n127) );
    zdffqrb DNT_DW10_Q_reg_31 ( .CK(DNT_DW10_n127), .D(ADI[31]), .R(TRST_), 
        .Q(DW10[31]) );
    zdffqrb DNT_DW10_Q_reg_30 ( .CK(DNT_DW10_n127), .D(ADI[30]), .R(TRST_), 
        .Q(DW10[30]) );
    zdffqrb DNT_DW10_Q_reg_29 ( .CK(DNT_DW10_n127), .D(ADI[29]), .R(TRST_), 
        .Q(DW10[29]) );
    zdffqrb DNT_DW10_Q_reg_28 ( .CK(DNT_DW10_n127), .D(ADI[28]), .R(TRST_), 
        .Q(DW10[28]) );
    zdffqrb DNT_DW10_Q_reg_27 ( .CK(DNT_DW10_n127), .D(ADI[27]), .R(TRST_), 
        .Q(DW10[27]) );
    zdffqrb DNT_DW10_Q_reg_26 ( .CK(DNT_DW10_n127), .D(ADI[26]), .R(TRST_), 
        .Q(DW10[26]) );
    zdffqrb DNT_DW10_Q_reg_25 ( .CK(DNT_DW10_n127), .D(ADI[25]), .R(TRST_), 
        .Q(DW10[25]) );
    zdffqrb DNT_DW10_Q_reg_24 ( .CK(DNT_DW10_n127), .D(ADI[24]), .R(TRST_), 
        .Q(DW10[24]) );
    zdffqrb DNT_DW10_Q_reg_23 ( .CK(DNT_DW10_n127), .D(ADI[23]), .R(TRST_), 
        .Q(DW10[23]) );
    zdffqrb DNT_DW10_Q_reg_22 ( .CK(DNT_DW10_n127), .D(ADI[22]), .R(TRST_), 
        .Q(DW10[22]) );
    zdffqrb DNT_DW10_Q_reg_21 ( .CK(DNT_DW10_n127), .D(ADI[21]), .R(TRST_), 
        .Q(DW10[21]) );
    zdffqrb DNT_DW10_Q_reg_20 ( .CK(DNT_DW10_n127), .D(ADI[20]), .R(TRST_), 
        .Q(DW10[20]) );
    zdffqrb DNT_DW10_Q_reg_19 ( .CK(DNT_DW10_n127), .D(ADI[19]), .R(TRST_), 
        .Q(DW10[19]) );
    zdffqrb DNT_DW10_Q_reg_18 ( .CK(DNT_DW10_n127), .D(ADI[18]), .R(TRST_), 
        .Q(DW10[18]) );
    zdffqrb DNT_DW10_Q_reg_17 ( .CK(DNT_DW10_n127), .D(ADI[17]), .R(TRST_), 
        .Q(DW10[17]) );
    zdffqrb DNT_DW10_Q_reg_16 ( .CK(DNT_DW10_n127), .D(ADI[16]), .R(TRST_), 
        .Q(DW10[16]) );
    zdffqrb DNT_DW10_Q_reg_15 ( .CK(DNT_DW10_n126), .D(ADI[15]), .R(TRST_), 
        .Q(DW10[15]) );
    zdffqrb DNT_DW10_Q_reg_14 ( .CK(DNT_DW10_n126), .D(ADI[14]), .R(TRST_), 
        .Q(DW10[14]) );
    zdffqrb DNT_DW10_Q_reg_13 ( .CK(DNT_DW10_n126), .D(ADI[13]), .R(TRST_), 
        .Q(DW10[13]) );
    zdffqrb DNT_DW10_Q_reg_12 ( .CK(DNT_DW10_n126), .D(ADI[12]), .R(TRST_), 
        .Q(DW10[12]) );
    zdffqrb DNT_DW10_Q_reg_11 ( .CK(DNT_DW10_n126), .D(ADI[11]), .R(TRST_), 
        .Q(DW10[11]) );
    zdffqrb DNT_DW10_Q_reg_10 ( .CK(DNT_DW10_n126), .D(ADI[10]), .R(TRST_), 
        .Q(DW10[10]) );
    zdffqrb DNT_DW10_Q_reg_9 ( .CK(DNT_DW10_n126), .D(ADI[9]), .R(TRST_), .Q(
        DW10[9]) );
    zdffqrb DNT_DW10_Q_reg_8 ( .CK(DNT_DW10_n126), .D(ADI[8]), .R(TRST_), .Q(
        DW10[8]) );
    zdffqrb DNT_DW10_Q_reg_7 ( .CK(DNT_DW10_n126), .D(ADI[7]), .R(TRST_), .Q(
        DW10[7]) );
    zdffqrb DNT_DW10_Q_reg_6 ( .CK(DNT_DW10_n126), .D(ADI[6]), .R(TRST_), .Q(
        DW10[6]) );
    zdffqrb DNT_DW10_Q_reg_5 ( .CK(DNT_DW10_n126), .D(ADI[5]), .R(TRST_), .Q(
        DW10[5]) );
    zdffqrb DNT_DW10_Q_reg_4 ( .CK(DNT_DW10_n126), .D(ADI[4]), .R(TRST_), .Q(
        DW10[4]) );
    zdffqrb DNT_DW10_Q_reg_3 ( .CK(DNT_DW10_n126), .D(ADI[3]), .R(TRST_), .Q(
        DW10[3]) );
    zdffqrb DNT_DW10_Q_reg_2 ( .CK(DNT_DW10_n126), .D(ADI[2]), .R(TRST_), .Q(
        DW10[2]) );
    zdffqrb DNT_DW10_Q_reg_1 ( .CK(DNT_DW10_n126), .D(ADI[1]), .R(TRST_), .Q(
        DW10[1]) );
    zdffqrb DNT_DW10_Q_reg_0 ( .CK(DNT_DW10_n126), .D(ADI[0]), .R(TRST_), .Q(
        DW10[0]) );
    zbfb DNT_DW10_U80 ( .A(FLOPS_CLK_14), .Y(DNT_DW10_n126) );
    zbfb DNT_DW10_U81 ( .A(FLOPS_CLK_14), .Y(DNT_DW10_n127) );
    zdffqrb DNT_DW8_Q_reg_31 ( .CK(DNT_DW8_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW8[31]) );
    zdffqrb DNT_DW8_Q_reg_30 ( .CK(DNT_DW8_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW8[30]) );
    zdffqrb DNT_DW8_Q_reg_29 ( .CK(DNT_DW8_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW8[29]) );
    zdffqrb DNT_DW8_Q_reg_28 ( .CK(DNT_DW8_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW8[28]) );
    zdffqrb DNT_DW8_Q_reg_27 ( .CK(DNT_DW8_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW8[27]) );
    zdffqrb DNT_DW8_Q_reg_26 ( .CK(DNT_DW8_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW8[26]) );
    zdffqrb DNT_DW8_Q_reg_25 ( .CK(DNT_DW8_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW8[25]) );
    zdffqrb DNT_DW8_Q_reg_24 ( .CK(DNT_DW8_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW8[24]) );
    zdffqrb DNT_DW8_Q_reg_23 ( .CK(DNT_DW8_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW8[23]) );
    zdffqrb DNT_DW8_Q_reg_22 ( .CK(DNT_DW8_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW8[22]) );
    zdffqrb DNT_DW8_Q_reg_21 ( .CK(DNT_DW8_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW8[21]) );
    zdffqrb DNT_DW8_Q_reg_20 ( .CK(DNT_DW8_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW8[20]) );
    zdffqrb DNT_DW8_Q_reg_19 ( .CK(DNT_DW8_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW8[19]) );
    zdffqrb DNT_DW8_Q_reg_18 ( .CK(DNT_DW8_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW8[18]) );
    zdffqrb DNT_DW8_Q_reg_17 ( .CK(DNT_DW8_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW8[17]) );
    zdffqrb DNT_DW8_Q_reg_16 ( .CK(DNT_DW8_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW8[16]) );
    zdffqrb DNT_DW8_Q_reg_15 ( .CK(DNT_DW8_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW8[15]) );
    zdffqrb DNT_DW8_Q_reg_14 ( .CK(DNT_DW8_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW8[14]) );
    zdffqrb DNT_DW8_Q_reg_13 ( .CK(DNT_DW8_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW8[13]) );
    zdffqrb DNT_DW8_Q_reg_12 ( .CK(DNT_DW8_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW8[12]) );
    zdffqrb DNT_DW8_Q_reg_11 ( .CK(DNT_DW8_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW8[11]) );
    zdffqrb DNT_DW8_Q_reg_10 ( .CK(DNT_DW8_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW8[10]) );
    zdffqrb DNT_DW8_Q_reg_9 ( .CK(DNT_DW8_n126), .D(ADI[9]), .R(TRST_), .Q(DW8
        [9]) );
    zdffqrb DNT_DW8_Q_reg_8 ( .CK(DNT_DW8_n126), .D(ADI[8]), .R(TRST_), .Q(DW8
        [8]) );
    zdffqrb DNT_DW8_Q_reg_7 ( .CK(DNT_DW8_n126), .D(ADI[7]), .R(TRST_), .Q(DW8
        [7]) );
    zdffqrb DNT_DW8_Q_reg_6 ( .CK(DNT_DW8_n126), .D(ADI[6]), .R(TRST_), .Q(DW8
        [6]) );
    zdffqrb DNT_DW8_Q_reg_5 ( .CK(DNT_DW8_n126), .D(ADI[5]), .R(TRST_), .Q(DW8
        [5]) );
    zdffqrb DNT_DW8_Q_reg_4 ( .CK(DNT_DW8_n126), .D(ADI[4]), .R(TRST_), .Q(DW8
        [4]) );
    zdffqrb DNT_DW8_Q_reg_3 ( .CK(DNT_DW8_n126), .D(ADI[3]), .R(TRST_), .Q(DW8
        [3]) );
    zdffqrb DNT_DW8_Q_reg_2 ( .CK(DNT_DW8_n126), .D(ADI[2]), .R(TRST_), .Q(DW8
        [2]) );
    zdffqrb DNT_DW8_Q_reg_1 ( .CK(DNT_DW8_n126), .D(ADI[1]), .R(TRST_), .Q(DW8
        [1]) );
    zdffqrb DNT_DW8_Q_reg_0 ( .CK(DNT_DW8_n126), .D(ADI[0]), .R(TRST_), .Q(DW8
        [0]) );
    zbfb DNT_DW8_U80 ( .A(FLOPS_CLK_12), .Y(DNT_DW8_n126) );
    zbfb DNT_DW8_U81 ( .A(FLOPS_CLK_12), .Y(DNT_DW8_n127) );
    zdffqrb DNT_DW0_Q_reg_31 ( .CK(DNT_DW0_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW0[31]) );
    zdffqrb DNT_DW0_Q_reg_30 ( .CK(DNT_DW0_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW0[30]) );
    zdffqrb DNT_DW0_Q_reg_29 ( .CK(DNT_DW0_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW0[29]) );
    zdffqrb DNT_DW0_Q_reg_28 ( .CK(DNT_DW0_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW0[28]) );
    zdffqrb DNT_DW0_Q_reg_27 ( .CK(DNT_DW0_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW0[27]) );
    zdffqrb DNT_DW0_Q_reg_26 ( .CK(DNT_DW0_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW0[26]) );
    zdffqrb DNT_DW0_Q_reg_25 ( .CK(DNT_DW0_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW0[25]) );
    zdffqrb DNT_DW0_Q_reg_24 ( .CK(DNT_DW0_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW0[24]) );
    zdffqrb DNT_DW0_Q_reg_23 ( .CK(DNT_DW0_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW0[23]) );
    zdffqrb DNT_DW0_Q_reg_22 ( .CK(DNT_DW0_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW0[22]) );
    zdffqrb DNT_DW0_Q_reg_21 ( .CK(DNT_DW0_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW0[21]) );
    zdffqrb DNT_DW0_Q_reg_20 ( .CK(DNT_DW0_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW0[20]) );
    zdffqrb DNT_DW0_Q_reg_19 ( .CK(DNT_DW0_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW0[19]) );
    zdffqrb DNT_DW0_Q_reg_18 ( .CK(DNT_DW0_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW0[18]) );
    zdffqrb DNT_DW0_Q_reg_17 ( .CK(DNT_DW0_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW0[17]) );
    zdffqrb DNT_DW0_Q_reg_16 ( .CK(DNT_DW0_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW0[16]) );
    zdffqrb DNT_DW0_Q_reg_15 ( .CK(DNT_DW0_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW0[15]) );
    zdffqrb DNT_DW0_Q_reg_14 ( .CK(DNT_DW0_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW0[14]) );
    zdffqrb DNT_DW0_Q_reg_13 ( .CK(DNT_DW0_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW0[13]) );
    zdffqrb DNT_DW0_Q_reg_12 ( .CK(DNT_DW0_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW0[12]) );
    zdffqrb DNT_DW0_Q_reg_11 ( .CK(DNT_DW0_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW0[11]) );
    zdffqrb DNT_DW0_Q_reg_10 ( .CK(DNT_DW0_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW0[10]) );
    zdffqrb DNT_DW0_Q_reg_9 ( .CK(DNT_DW0_n126), .D(ADI[9]), .R(TRST_), .Q(DW0
        [9]) );
    zdffqrb DNT_DW0_Q_reg_8 ( .CK(DNT_DW0_n126), .D(ADI[8]), .R(TRST_), .Q(DW0
        [8]) );
    zdffqrb DNT_DW0_Q_reg_7 ( .CK(DNT_DW0_n126), .D(ADI[7]), .R(TRST_), .Q(DW0
        [7]) );
    zdffqrb DNT_DW0_Q_reg_6 ( .CK(DNT_DW0_n126), .D(ADI[6]), .R(TRST_), .Q(DW0
        [6]) );
    zdffqrb DNT_DW0_Q_reg_5 ( .CK(DNT_DW0_n126), .D(ADI[5]), .R(TRST_), .Q(DW0
        [5]) );
    zdffqrb DNT_DW0_Q_reg_4 ( .CK(DNT_DW0_n126), .D(ADI[4]), .R(TRST_), .Q(DW0
        [4]) );
    zdffqrb DNT_DW0_Q_reg_3 ( .CK(DNT_DW0_n126), .D(ADI[3]), .R(TRST_), .Q(DW0
        [3]) );
    zdffqrb DNT_DW0_Q_reg_2 ( .CK(DNT_DW0_n126), .D(ADI[2]), .R(TRST_), .Q(DW0
        [2]) );
    zdffqrb DNT_DW0_Q_reg_1 ( .CK(DNT_DW0_n126), .D(ADI[1]), .R(TRST_), .Q(DW0
        [1]) );
    zdffqrb DNT_DW0_Q_reg_0 ( .CK(DNT_DW0_n126), .D(ADI[0]), .R(TRST_), .Q(DW0
        [0]) );
    zbfb DNT_DW0_U80 ( .A(FLOPS_CLK_4), .Y(DNT_DW0_n126) );
    zbfb DNT_DW0_U81 ( .A(FLOPS_CLK_4), .Y(DNT_DW0_n127) );
    zdffqrb DNT_DW11_Q_reg_31 ( .CK(DNT_DW11_n127), .D(ADI[31]), .R(TRST_), 
        .Q(DW11[31]) );
    zdffqrb DNT_DW11_Q_reg_30 ( .CK(DNT_DW11_n127), .D(ADI[30]), .R(TRST_), 
        .Q(DW11[30]) );
    zdffqrb DNT_DW11_Q_reg_29 ( .CK(DNT_DW11_n127), .D(ADI[29]), .R(TRST_), 
        .Q(DW11[29]) );
    zdffqrb DNT_DW11_Q_reg_28 ( .CK(DNT_DW11_n127), .D(ADI[28]), .R(TRST_), 
        .Q(DW11[28]) );
    zdffqrb DNT_DW11_Q_reg_27 ( .CK(DNT_DW11_n127), .D(ADI[27]), .R(TRST_), 
        .Q(DW11[27]) );
    zdffqrb DNT_DW11_Q_reg_26 ( .CK(DNT_DW11_n127), .D(ADI[26]), .R(TRST_), 
        .Q(DW11[26]) );
    zdffqrb DNT_DW11_Q_reg_25 ( .CK(DNT_DW11_n127), .D(ADI[25]), .R(TRST_), 
        .Q(DW11[25]) );
    zdffqrb DNT_DW11_Q_reg_24 ( .CK(DNT_DW11_n127), .D(ADI[24]), .R(TRST_), 
        .Q(DW11[24]) );
    zdffqrb DNT_DW11_Q_reg_23 ( .CK(DNT_DW11_n127), .D(ADI[23]), .R(TRST_), 
        .Q(DW11[23]) );
    zdffqrb DNT_DW11_Q_reg_22 ( .CK(DNT_DW11_n127), .D(ADI[22]), .R(TRST_), 
        .Q(DW11[22]) );
    zdffqrb DNT_DW11_Q_reg_21 ( .CK(DNT_DW11_n127), .D(ADI[21]), .R(TRST_), 
        .Q(DW11[21]) );
    zdffqrb DNT_DW11_Q_reg_20 ( .CK(DNT_DW11_n127), .D(ADI[20]), .R(TRST_), 
        .Q(DW11[20]) );
    zdffqrb DNT_DW11_Q_reg_19 ( .CK(DNT_DW11_n127), .D(ADI[19]), .R(TRST_), 
        .Q(DW11[19]) );
    zdffqrb DNT_DW11_Q_reg_18 ( .CK(DNT_DW11_n127), .D(ADI[18]), .R(TRST_), 
        .Q(DW11[18]) );
    zdffqrb DNT_DW11_Q_reg_17 ( .CK(DNT_DW11_n127), .D(ADI[17]), .R(TRST_), 
        .Q(DW11[17]) );
    zdffqrb DNT_DW11_Q_reg_16 ( .CK(DNT_DW11_n127), .D(ADI[16]), .R(TRST_), 
        .Q(DW11[16]) );
    zdffqrb DNT_DW11_Q_reg_15 ( .CK(DNT_DW11_n126), .D(ADI[15]), .R(TRST_), 
        .Q(DW11[15]) );
    zdffqrb DNT_DW11_Q_reg_14 ( .CK(DNT_DW11_n126), .D(ADI[14]), .R(TRST_), 
        .Q(DW11[14]) );
    zdffqrb DNT_DW11_Q_reg_13 ( .CK(DNT_DW11_n126), .D(ADI[13]), .R(TRST_), 
        .Q(DW11[13]) );
    zdffqrb DNT_DW11_Q_reg_12 ( .CK(DNT_DW11_n126), .D(ADI[12]), .R(TRST_), 
        .Q(DW11[12]) );
    zdffqrb DNT_DW11_Q_reg_11 ( .CK(DNT_DW11_n126), .D(ADI[11]), .R(TRST_), 
        .Q(DW11[11]) );
    zdffqrb DNT_DW11_Q_reg_10 ( .CK(DNT_DW11_n126), .D(ADI[10]), .R(TRST_), 
        .Q(DW11[10]) );
    zdffqrb DNT_DW11_Q_reg_9 ( .CK(DNT_DW11_n126), .D(ADI[9]), .R(TRST_), .Q(
        DW11[9]) );
    zdffqrb DNT_DW11_Q_reg_8 ( .CK(DNT_DW11_n126), .D(ADI[8]), .R(TRST_), .Q(
        DW11[8]) );
    zdffqrb DNT_DW11_Q_reg_7 ( .CK(DNT_DW11_n126), .D(ADI[7]), .R(TRST_), .Q(
        DW11[7]) );
    zdffqrb DNT_DW11_Q_reg_6 ( .CK(DNT_DW11_n126), .D(ADI[6]), .R(TRST_), .Q(
        DW11[6]) );
    zdffqrb DNT_DW11_Q_reg_5 ( .CK(DNT_DW11_n126), .D(ADI[5]), .R(TRST_), .Q(
        DW11[5]) );
    zdffqrb DNT_DW11_Q_reg_4 ( .CK(DNT_DW11_n126), .D(ADI[4]), .R(TRST_), .Q(
        DW11[4]) );
    zdffqrb DNT_DW11_Q_reg_3 ( .CK(DNT_DW11_n126), .D(ADI[3]), .R(TRST_), .Q(
        DW11[3]) );
    zdffqrb DNT_DW11_Q_reg_2 ( .CK(DNT_DW11_n126), .D(ADI[2]), .R(TRST_), .Q(
        DW11[2]) );
    zdffqrb DNT_DW11_Q_reg_1 ( .CK(DNT_DW11_n126), .D(ADI[1]), .R(TRST_), .Q(
        DW11[1]) );
    zdffqrb DNT_DW11_Q_reg_0 ( .CK(DNT_DW11_n126), .D(ADI[0]), .R(TRST_), .Q(
        DW11[0]) );
    zbfb DNT_DW11_U80 ( .A(FLOPS_CLK_15), .Y(DNT_DW11_n126) );
    zbfb DNT_DW11_U81 ( .A(FLOPS_CLK_15), .Y(DNT_DW11_n127) );
    zdffqrb DNT_DW9_Q_reg_31 ( .CK(DNT_DW9_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW9[31]) );
    zdffqrb DNT_DW9_Q_reg_30 ( .CK(DNT_DW9_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW9[30]) );
    zdffqrb DNT_DW9_Q_reg_29 ( .CK(DNT_DW9_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW9[29]) );
    zdffqrb DNT_DW9_Q_reg_28 ( .CK(DNT_DW9_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW9[28]) );
    zdffqrb DNT_DW9_Q_reg_27 ( .CK(DNT_DW9_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW9[27]) );
    zdffqrb DNT_DW9_Q_reg_26 ( .CK(DNT_DW9_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW9[26]) );
    zdffqrb DNT_DW9_Q_reg_25 ( .CK(DNT_DW9_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW9[25]) );
    zdffqrb DNT_DW9_Q_reg_24 ( .CK(DNT_DW9_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW9[24]) );
    zdffqrb DNT_DW9_Q_reg_23 ( .CK(DNT_DW9_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW9[23]) );
    zdffqrb DNT_DW9_Q_reg_22 ( .CK(DNT_DW9_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW9[22]) );
    zdffqrb DNT_DW9_Q_reg_21 ( .CK(DNT_DW9_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW9[21]) );
    zdffqrb DNT_DW9_Q_reg_20 ( .CK(DNT_DW9_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW9[20]) );
    zdffqrb DNT_DW9_Q_reg_19 ( .CK(DNT_DW9_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW9[19]) );
    zdffqrb DNT_DW9_Q_reg_18 ( .CK(DNT_DW9_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW9[18]) );
    zdffqrb DNT_DW9_Q_reg_17 ( .CK(DNT_DW9_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW9[17]) );
    zdffqrb DNT_DW9_Q_reg_16 ( .CK(DNT_DW9_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW9[16]) );
    zdffqrb DNT_DW9_Q_reg_15 ( .CK(DNT_DW9_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW9[15]) );
    zdffqrb DNT_DW9_Q_reg_14 ( .CK(DNT_DW9_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW9[14]) );
    zdffqrb DNT_DW9_Q_reg_13 ( .CK(DNT_DW9_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW9[13]) );
    zdffqrb DNT_DW9_Q_reg_12 ( .CK(DNT_DW9_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW9[12]) );
    zdffqrb DNT_DW9_Q_reg_11 ( .CK(DNT_DW9_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW9[11]) );
    zdffqrb DNT_DW9_Q_reg_10 ( .CK(DNT_DW9_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW9[10]) );
    zdffqrb DNT_DW9_Q_reg_9 ( .CK(DNT_DW9_n126), .D(ADI[9]), .R(TRST_), .Q(DW9
        [9]) );
    zdffqrb DNT_DW9_Q_reg_8 ( .CK(DNT_DW9_n126), .D(ADI[8]), .R(TRST_), .Q(DW9
        [8]) );
    zdffqrb DNT_DW9_Q_reg_7 ( .CK(DNT_DW9_n126), .D(ADI[7]), .R(TRST_), .Q(DW9
        [7]) );
    zdffqrb DNT_DW9_Q_reg_6 ( .CK(DNT_DW9_n126), .D(ADI[6]), .R(TRST_), .Q(DW9
        [6]) );
    zdffqrb DNT_DW9_Q_reg_5 ( .CK(DNT_DW9_n126), .D(ADI[5]), .R(TRST_), .Q(DW9
        [5]) );
    zdffqrb DNT_DW9_Q_reg_4 ( .CK(DNT_DW9_n126), .D(ADI[4]), .R(TRST_), .Q(DW9
        [4]) );
    zdffqrb DNT_DW9_Q_reg_3 ( .CK(DNT_DW9_n126), .D(ADI[3]), .R(TRST_), .Q(DW9
        [3]) );
    zdffqrb DNT_DW9_Q_reg_2 ( .CK(DNT_DW9_n126), .D(ADI[2]), .R(TRST_), .Q(DW9
        [2]) );
    zdffqrb DNT_DW9_Q_reg_1 ( .CK(DNT_DW9_n126), .D(ADI[1]), .R(TRST_), .Q(DW9
        [1]) );
    zdffqrb DNT_DW9_Q_reg_0 ( .CK(DNT_DW9_n126), .D(ADI[0]), .R(TRST_), .Q(DW9
        [0]) );
    zbfb DNT_DW9_U80 ( .A(FLOPS_CLK_13), .Y(DNT_DW9_n126) );
    zbfb DNT_DW9_U81 ( .A(FLOPS_CLK_13), .Y(DNT_DW9_n127) );
    zdffqrb DNT_DW7_Q_reg_31 ( .CK(DNT_DW7_n127), .D(AD7IN_31), .R(TRST_), .Q(
        DW7[31]) );
    zdffqrb DNT_DW7_Q_reg_30 ( .CK(DNT_DW7_n127), .D(AD7IN_30), .R(TRST_), .Q(
        DW7[30]) );
    zdffqrb DNT_DW7_Q_reg_29 ( .CK(DNT_DW7_n127), .D(AD7IN_29), .R(TRST_), .Q(
        DW7[29]) );
    zdffqrb DNT_DW7_Q_reg_28 ( .CK(DNT_DW7_n127), .D(AD7IN_28), .R(TRST_), .Q(
        DW7[28]) );
    zdffqrb DNT_DW7_Q_reg_27 ( .CK(DNT_DW7_n127), .D(AD7IN_27), .R(TRST_), .Q(
        DW7[27]) );
    zdffqrb DNT_DW7_Q_reg_26 ( .CK(DNT_DW7_n127), .D(AD7IN_26), .R(TRST_), .Q(
        DW7[26]) );
    zdffqrb DNT_DW7_Q_reg_25 ( .CK(DNT_DW7_n127), .D(AD7IN_25), .R(TRST_), .Q(
        DW7[25]) );
    zdffqrb DNT_DW7_Q_reg_24 ( .CK(DNT_DW7_n127), .D(AD7IN_24), .R(TRST_), .Q(
        DW7[24]) );
    zdffqrb DNT_DW7_Q_reg_23 ( .CK(DNT_DW7_n127), .D(AD7IN_23), .R(TRST_), .Q(
        DW7[23]) );
    zdffqrb DNT_DW7_Q_reg_22 ( .CK(DNT_DW7_n127), .D(AD7IN_22), .R(TRST_), .Q(
        DW7[22]) );
    zdffqrb DNT_DW7_Q_reg_21 ( .CK(DNT_DW7_n127), .D(AD7IN_21), .R(TRST_), .Q(
        DW7[21]) );
    zdffqrb DNT_DW7_Q_reg_20 ( .CK(DNT_DW7_n127), .D(AD7IN_20), .R(TRST_), .Q(
        DW7[20]) );
    zdffqrb DNT_DW7_Q_reg_19 ( .CK(DNT_DW7_n127), .D(AD7IN_19), .R(TRST_), .Q(
        DW7[19]) );
    zdffqrb DNT_DW7_Q_reg_18 ( .CK(DNT_DW7_n127), .D(AD7IN_18), .R(TRST_), .Q(
        DW7[18]) );
    zdffqrb DNT_DW7_Q_reg_17 ( .CK(DNT_DW7_n127), .D(AD7IN_17), .R(TRST_), .Q(
        DW7[17]) );
    zdffqrb DNT_DW7_Q_reg_16 ( .CK(DNT_DW7_n127), .D(AD7IN_16), .R(TRST_), .Q(
        DW7[16]) );
    zdffqrb DNT_DW7_Q_reg_15 ( .CK(DNT_DW7_n126), .D(AD7IN_15), .R(TRST_), .Q(
        DW7[15]) );
    zdffqrb DNT_DW7_Q_reg_14 ( .CK(DNT_DW7_n126), .D(AD7IN_14), .R(TRST_), .Q(
        DW7[14]) );
    zdffqrb DNT_DW7_Q_reg_13 ( .CK(DNT_DW7_n126), .D(AD7IN_13), .R(TRST_), .Q(
        DW7[13]) );
    zdffqrb DNT_DW7_Q_reg_12 ( .CK(DNT_DW7_n126), .D(AD7IN_12), .R(TRST_), .Q(
        DW7[12]) );
    zdffqrb DNT_DW7_Q_reg_11 ( .CK(DNT_DW7_n126), .D(AD7IN_11), .R(TRST_), .Q(
        DW7[11]) );
    zdffqrb DNT_DW7_Q_reg_10 ( .CK(DNT_DW7_n126), .D(AD7IN_10), .R(TRST_), .Q(
        DW7[10]) );
    zdffqrb DNT_DW7_Q_reg_9 ( .CK(DNT_DW7_n126), .D(AD7IN_9), .R(TRST_), .Q(
        DW7[9]) );
    zdffqrb DNT_DW7_Q_reg_8 ( .CK(DNT_DW7_n126), .D(AD7IN_8), .R(TRST_), .Q(
        DW7[8]) );
    zdffqrb DNT_DW7_Q_reg_7 ( .CK(DNT_DW7_n126), .D(AD7IN_7), .R(TRST_), .Q(
        DW7[7]) );
    zdffqrb DNT_DW7_Q_reg_6 ( .CK(DNT_DW7_n126), .D(AD7IN_6), .R(TRST_), .Q(
        DW7[6]) );
    zdffqrb DNT_DW7_Q_reg_5 ( .CK(DNT_DW7_n126), .D(AD7IN_5), .R(TRST_), .Q(
        DW7[5]) );
    zdffqrb DNT_DW7_Q_reg_4 ( .CK(DNT_DW7_n126), .D(AD7IN_4), .R(TRST_), .Q(
        DW7[4]) );
    zdffqrb DNT_DW7_Q_reg_3 ( .CK(DNT_DW7_n126), .D(AD7IN_3), .R(TRST_), .Q(
        DW7[3]) );
    zdffqrb DNT_DW7_Q_reg_2 ( .CK(DNT_DW7_n126), .D(AD7IN_2), .R(TRST_), .Q(
        DW7[2]) );
    zdffqrb DNT_DW7_Q_reg_1 ( .CK(DNT_DW7_n126), .D(AD7IN_1), .R(TRST_), .Q(
        DW7[1]) );
    zdffqrb DNT_DW7_Q_reg_0 ( .CK(DNT_DW7_n126), .D(AD7IN_0), .R(TRST_), .Q(
        DW7[0]) );
    zbfb DNT_DW7_U80 ( .A(FLOPS_CLK_11), .Y(DNT_DW7_n126) );
    zbfb DNT_DW7_U81 ( .A(FLOPS_CLK_11), .Y(DNT_DW7_n127) );
    zdffqrb DNT_DW5_Q_reg_31 ( .CK(DNT_DW5_n127), .D(AD5IN_31), .R(TRST_), .Q(
        DW5[31]) );
    zdffqrb DNT_DW5_Q_reg_30 ( .CK(DNT_DW5_n127), .D(AD5IN_30), .R(TRST_), .Q(
        DW5[30]) );
    zdffqrb DNT_DW5_Q_reg_29 ( .CK(DNT_DW5_n127), .D(AD5IN_29), .R(TRST_), .Q(
        DW5[29]) );
    zdffqrb DNT_DW5_Q_reg_28 ( .CK(DNT_DW5_n127), .D(AD5IN_28), .R(TRST_), .Q(
        DW5[28]) );
    zdffqrb DNT_DW5_Q_reg_27 ( .CK(DNT_DW5_n127), .D(AD5IN_27), .R(TRST_), .Q(
        DW5[27]) );
    zdffqrb DNT_DW5_Q_reg_26 ( .CK(DNT_DW5_n127), .D(AD5IN_26), .R(TRST_), .Q(
        DW5[26]) );
    zdffqrb DNT_DW5_Q_reg_25 ( .CK(DNT_DW5_n127), .D(AD5IN_25), .R(TRST_), .Q(
        DW5[25]) );
    zdffqrb DNT_DW5_Q_reg_24 ( .CK(DNT_DW5_n127), .D(AD5IN_24), .R(TRST_), .Q(
        DW5[24]) );
    zdffqrb DNT_DW5_Q_reg_23 ( .CK(DNT_DW5_n127), .D(AD5IN_23), .R(TRST_), .Q(
        DW5[23]) );
    zdffqrb DNT_DW5_Q_reg_22 ( .CK(DNT_DW5_n127), .D(AD5IN_22), .R(TRST_), .Q(
        DW5[22]) );
    zdffqrb DNT_DW5_Q_reg_21 ( .CK(DNT_DW5_n127), .D(AD5IN_21), .R(TRST_), .Q(
        DW5[21]) );
    zdffqrb DNT_DW5_Q_reg_20 ( .CK(DNT_DW5_n127), .D(AD5IN_20), .R(TRST_), .Q(
        DW5[20]) );
    zdffqrb DNT_DW5_Q_reg_19 ( .CK(DNT_DW5_n127), .D(AD5IN_19), .R(TRST_), .Q(
        DW5[19]) );
    zdffqrb DNT_DW5_Q_reg_18 ( .CK(DNT_DW5_n127), .D(AD5IN_18), .R(TRST_), .Q(
        DW5[18]) );
    zdffqrb DNT_DW5_Q_reg_17 ( .CK(DNT_DW5_n127), .D(AD5IN_17), .R(TRST_), .Q(
        DW5[17]) );
    zdffqrb DNT_DW5_Q_reg_16 ( .CK(DNT_DW5_n127), .D(AD5IN_16), .R(TRST_), .Q(
        DW5[16]) );
    zdffqrb DNT_DW5_Q_reg_15 ( .CK(DNT_DW5_n126), .D(AD5IN_15), .R(TRST_), .Q(
        DW5[15]) );
    zdffqrb DNT_DW5_Q_reg_14 ( .CK(DNT_DW5_n126), .D(AD5IN_14), .R(TRST_), .Q(
        DW5[14]) );
    zdffqrb DNT_DW5_Q_reg_13 ( .CK(DNT_DW5_n126), .D(AD5IN_13), .R(TRST_), .Q(
        DW5[13]) );
    zdffqrb DNT_DW5_Q_reg_12 ( .CK(DNT_DW5_n126), .D(AD5IN_12), .R(TRST_), .Q(
        DW5[12]) );
    zdffqrb DNT_DW5_Q_reg_11 ( .CK(DNT_DW5_n126), .D(AD5IN_11), .R(TRST_), .Q(
        DW5[11]) );
    zdffqrb DNT_DW5_Q_reg_10 ( .CK(DNT_DW5_n126), .D(AD5IN_10), .R(TRST_), .Q(
        DW5[10]) );
    zdffqrb DNT_DW5_Q_reg_9 ( .CK(DNT_DW5_n126), .D(AD5IN_9), .R(TRST_), .Q(
        DW5[9]) );
    zdffqrb DNT_DW5_Q_reg_8 ( .CK(DNT_DW5_n126), .D(AD5IN_8), .R(TRST_), .Q(
        DW5[8]) );
    zdffqrb DNT_DW5_Q_reg_7 ( .CK(DNT_DW5_n126), .D(AD5IN_7), .R(TRST_), .Q(
        DW5[7]) );
    zdffqrb DNT_DW5_Q_reg_6 ( .CK(DNT_DW5_n126), .D(AD5IN_6), .R(TRST_), .Q(
        DW5[6]) );
    zdffqrb DNT_DW5_Q_reg_5 ( .CK(DNT_DW5_n126), .D(AD5IN_5), .R(TRST_), .Q(
        DW5[5]) );
    zdffqrb DNT_DW5_Q_reg_4 ( .CK(DNT_DW5_n126), .D(AD5IN_4), .R(TRST_), .Q(
        DW5[4]) );
    zdffqrb DNT_DW5_Q_reg_3 ( .CK(DNT_DW5_n126), .D(AD5IN_3), .R(TRST_), .Q(
        DW5[3]) );
    zdffqrb DNT_DW5_Q_reg_2 ( .CK(DNT_DW5_n126), .D(AD5IN_2), .R(TRST_), .Q(
        DW5[2]) );
    zdffqrb DNT_DW5_Q_reg_1 ( .CK(DNT_DW5_n126), .D(AD5IN_1), .R(TRST_), .Q(
        DW5[1]) );
    zdffqrb DNT_DW5_Q_reg_0 ( .CK(DNT_DW5_n126), .D(AD5IN_0), .R(TRST_), .Q(
        DW5[0]) );
    zbfb DNT_DW5_U80 ( .A(FLOPS_CLK_9), .Y(DNT_DW5_n126) );
    zbfb DNT_DW5_U81 ( .A(FLOPS_CLK_9), .Y(DNT_DW5_n127) );
    zdffqrb DNT_DW2_Q_reg_31 ( .CK(DNT_DW2_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW2[31]) );
    zdffqrb DNT_DW2_Q_reg_30 ( .CK(DNT_DW2_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW2[30]) );
    zdffqrb DNT_DW2_Q_reg_29 ( .CK(DNT_DW2_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW2[29]) );
    zdffqrb DNT_DW2_Q_reg_28 ( .CK(DNT_DW2_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW2[28]) );
    zdffqrb DNT_DW2_Q_reg_27 ( .CK(DNT_DW2_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW2[27]) );
    zdffqrb DNT_DW2_Q_reg_26 ( .CK(DNT_DW2_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW2[26]) );
    zdffqrb DNT_DW2_Q_reg_25 ( .CK(DNT_DW2_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW2[25]) );
    zdffqrb DNT_DW2_Q_reg_24 ( .CK(DNT_DW2_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW2[24]) );
    zdffqrb DNT_DW2_Q_reg_23 ( .CK(DNT_DW2_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW2[23]) );
    zdffqrb DNT_DW2_Q_reg_22 ( .CK(DNT_DW2_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW2[22]) );
    zdffqrb DNT_DW2_Q_reg_21 ( .CK(DNT_DW2_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW2[21]) );
    zdffqrb DNT_DW2_Q_reg_20 ( .CK(DNT_DW2_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW2[20]) );
    zdffqrb DNT_DW2_Q_reg_19 ( .CK(DNT_DW2_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW2[19]) );
    zdffqrb DNT_DW2_Q_reg_18 ( .CK(DNT_DW2_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW2[18]) );
    zdffqrb DNT_DW2_Q_reg_17 ( .CK(DNT_DW2_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW2[17]) );
    zdffqrb DNT_DW2_Q_reg_16 ( .CK(DNT_DW2_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW2[16]) );
    zdffqrb DNT_DW2_Q_reg_15 ( .CK(DNT_DW2_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW2[15]) );
    zdffqrb DNT_DW2_Q_reg_14 ( .CK(DNT_DW2_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW2[14]) );
    zdffqrb DNT_DW2_Q_reg_13 ( .CK(DNT_DW2_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW2[13]) );
    zdffqrb DNT_DW2_Q_reg_12 ( .CK(DNT_DW2_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW2[12]) );
    zdffqrb DNT_DW2_Q_reg_11 ( .CK(DNT_DW2_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW2[11]) );
    zdffqrb DNT_DW2_Q_reg_10 ( .CK(DNT_DW2_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW2[10]) );
    zdffqrb DNT_DW2_Q_reg_9 ( .CK(DNT_DW2_n126), .D(ADI[9]), .R(TRST_), .Q(DW2
        [9]) );
    zdffqrb DNT_DW2_Q_reg_8 ( .CK(DNT_DW2_n126), .D(ADI[8]), .R(TRST_), .Q(DW2
        [8]) );
    zdffqrb DNT_DW2_Q_reg_7 ( .CK(DNT_DW2_n126), .D(ADI[7]), .R(TRST_), .Q(DW2
        [7]) );
    zdffqrb DNT_DW2_Q_reg_6 ( .CK(DNT_DW2_n126), .D(ADI[6]), .R(TRST_), .Q(DW2
        [6]) );
    zdffqrb DNT_DW2_Q_reg_5 ( .CK(DNT_DW2_n126), .D(ADI[5]), .R(TRST_), .Q(DW2
        [5]) );
    zdffqrb DNT_DW2_Q_reg_4 ( .CK(DNT_DW2_n126), .D(ADI[4]), .R(TRST_), .Q(DW2
        [4]) );
    zdffqrb DNT_DW2_Q_reg_3 ( .CK(DNT_DW2_n126), .D(ADI[3]), .R(TRST_), .Q(DW2
        [3]) );
    zdffqrb DNT_DW2_Q_reg_2 ( .CK(DNT_DW2_n126), .D(ADI[2]), .R(TRST_), .Q(DW2
        [2]) );
    zdffqrb DNT_DW2_Q_reg_1 ( .CK(DNT_DW2_n126), .D(ADI[1]), .R(TRST_), .Q(DW2
        [1]) );
    zdffqrb DNT_DW2_Q_reg_0 ( .CK(DNT_DW2_n126), .D(ADI[0]), .R(TRST_), .Q(DW2
        [0]) );
    zbfb DNT_DW2_U80 ( .A(FLOPS_CLK_6), .Y(DNT_DW2_n126) );
    zbfb DNT_DW2_U81 ( .A(FLOPS_CLK_6), .Y(DNT_DW2_n127) );
    zdffqrb DNT_DW3_Q_reg_31 ( .CK(DNT_DW3_n127), .D(AD3IN_31), .R(TRST_), .Q(
        DW3[31]) );
    zdffqrb DNT_DW3_Q_reg_30 ( .CK(DNT_DW3_n127), .D(AD3IN_30), .R(TRST_), .Q(
        DW3[30]) );
    zdffqrb DNT_DW3_Q_reg_29 ( .CK(DNT_DW3_n127), .D(AD3IN_29), .R(TRST_), .Q(
        DW3[29]) );
    zdffqrb DNT_DW3_Q_reg_28 ( .CK(DNT_DW3_n127), .D(AD3IN_28), .R(TRST_), .Q(
        DW3[28]) );
    zdffqrb DNT_DW3_Q_reg_27 ( .CK(DNT_DW3_n127), .D(AD3IN_27), .R(TRST_), .Q(
        DW3[27]) );
    zdffqrb DNT_DW3_Q_reg_26 ( .CK(DNT_DW3_n127), .D(AD3IN_26), .R(TRST_), .Q(
        DW3[26]) );
    zdffqrb DNT_DW3_Q_reg_25 ( .CK(DNT_DW3_n127), .D(AD3IN_25), .R(TRST_), .Q(
        DW3[25]) );
    zdffqrb DNT_DW3_Q_reg_24 ( .CK(DNT_DW3_n127), .D(AD3IN_24), .R(TRST_), .Q(
        DW3[24]) );
    zdffqrb DNT_DW3_Q_reg_23 ( .CK(DNT_DW3_n127), .D(AD3IN_23), .R(TRST_), .Q(
        DW3[23]) );
    zdffqrb DNT_DW3_Q_reg_22 ( .CK(DNT_DW3_n127), .D(AD3IN_22), .R(TRST_), .Q(
        DW3[22]) );
    zdffqrb DNT_DW3_Q_reg_21 ( .CK(DNT_DW3_n127), .D(AD3IN_21), .R(TRST_), .Q(
        DW3[21]) );
    zdffqrb DNT_DW3_Q_reg_20 ( .CK(DNT_DW3_n127), .D(AD3IN_20), .R(TRST_), .Q(
        DW3[20]) );
    zdffqrb DNT_DW3_Q_reg_19 ( .CK(DNT_DW3_n127), .D(AD3IN_19), .R(TRST_), .Q(
        DW3[19]) );
    zdffqrb DNT_DW3_Q_reg_18 ( .CK(DNT_DW3_n127), .D(AD3IN_18), .R(TRST_), .Q(
        DW3[18]) );
    zdffqrb DNT_DW3_Q_reg_17 ( .CK(DNT_DW3_n127), .D(AD3IN_17), .R(TRST_), .Q(
        DW3[17]) );
    zdffqrb DNT_DW3_Q_reg_16 ( .CK(DNT_DW3_n127), .D(AD3IN_16), .R(TRST_), .Q(
        DW3[16]) );
    zdffqrb DNT_DW3_Q_reg_15 ( .CK(DNT_DW3_n126), .D(AD3IN_15), .R(TRST_), .Q(
        DW3[15]) );
    zdffqrb DNT_DW3_Q_reg_14 ( .CK(DNT_DW3_n126), .D(AD3IN_14), .R(TRST_), .Q(
        DW3[14]) );
    zdffqrb DNT_DW3_Q_reg_13 ( .CK(DNT_DW3_n126), .D(AD3IN_13), .R(TRST_), .Q(
        DW3[13]) );
    zdffqrb DNT_DW3_Q_reg_12 ( .CK(DNT_DW3_n126), .D(AD3IN_12), .R(TRST_), .Q(
        DW3[12]) );
    zdffqrb DNT_DW3_Q_reg_11 ( .CK(DNT_DW3_n126), .D(AD3IN_11), .R(TRST_), .Q(
        DW3[11]) );
    zdffqrb DNT_DW3_Q_reg_10 ( .CK(DNT_DW3_n126), .D(AD3IN_10), .R(TRST_), .Q(
        DW3[10]) );
    zdffqrb DNT_DW3_Q_reg_9 ( .CK(DNT_DW3_n126), .D(AD3IN_9), .R(TRST_), .Q(
        DW3[9]) );
    zdffqrb DNT_DW3_Q_reg_8 ( .CK(DNT_DW3_n126), .D(AD3IN_8), .R(TRST_), .Q(
        DW3[8]) );
    zdffqrb DNT_DW3_Q_reg_7 ( .CK(DNT_DW3_n126), .D(AD3IN_7), .R(TRST_), .Q(
        DW3[7]) );
    zdffqrb DNT_DW3_Q_reg_6 ( .CK(DNT_DW3_n126), .D(AD3IN_6), .R(TRST_), .Q(
        DW3[6]) );
    zdffqrb DNT_DW3_Q_reg_5 ( .CK(DNT_DW3_n126), .D(AD3IN_5), .R(TRST_), .Q(
        DW3[5]) );
    zdffqrb DNT_DW3_Q_reg_4 ( .CK(DNT_DW3_n126), .D(AD3IN_4), .R(TRST_), .Q(
        DW3[4]) );
    zdffqrb DNT_DW3_Q_reg_3 ( .CK(DNT_DW3_n126), .D(AD3IN_3), .R(TRST_), .Q(
        DW3[3]) );
    zdffqrb DNT_DW3_Q_reg_2 ( .CK(DNT_DW3_n126), .D(AD3IN_2), .R(TRST_), .Q(
        DW3[2]) );
    zdffqrb DNT_DW3_Q_reg_1 ( .CK(DNT_DW3_n126), .D(AD3IN_1), .R(TRST_), .Q(
        DW3[1]) );
    zdffqrb DNT_DW3_Q_reg_0 ( .CK(DNT_DW3_n126), .D(AD3IN_0), .R(TRST_), .Q(
        DW3[0]) );
    zbfb DNT_DW3_U80 ( .A(FLOPS_CLK_7), .Y(DNT_DW3_n126) );
    zbfb DNT_DW3_U81 ( .A(FLOPS_CLK_7), .Y(DNT_DW3_n127) );
    zdffqrb DNT_DW4_Q_reg_31 ( .CK(DNT_DW4_n127), .D(ADI[31]), .R(TRST_), .Q(
        DW4[31]) );
    zdffqrb DNT_DW4_Q_reg_30 ( .CK(DNT_DW4_n127), .D(ADI[30]), .R(TRST_), .Q(
        DW4[30]) );
    zdffqrb DNT_DW4_Q_reg_29 ( .CK(DNT_DW4_n127), .D(ADI[29]), .R(TRST_), .Q(
        DW4[29]) );
    zdffqrb DNT_DW4_Q_reg_28 ( .CK(DNT_DW4_n127), .D(ADI[28]), .R(TRST_), .Q(
        DW4[28]) );
    zdffqrb DNT_DW4_Q_reg_27 ( .CK(DNT_DW4_n127), .D(ADI[27]), .R(TRST_), .Q(
        DW4[27]) );
    zdffqrb DNT_DW4_Q_reg_26 ( .CK(DNT_DW4_n127), .D(ADI[26]), .R(TRST_), .Q(
        DW4[26]) );
    zdffqrb DNT_DW4_Q_reg_25 ( .CK(DNT_DW4_n127), .D(ADI[25]), .R(TRST_), .Q(
        DW4[25]) );
    zdffqrb DNT_DW4_Q_reg_24 ( .CK(DNT_DW4_n127), .D(ADI[24]), .R(TRST_), .Q(
        DW4[24]) );
    zdffqrb DNT_DW4_Q_reg_23 ( .CK(DNT_DW4_n127), .D(ADI[23]), .R(TRST_), .Q(
        DW4[23]) );
    zdffqrb DNT_DW4_Q_reg_22 ( .CK(DNT_DW4_n127), .D(ADI[22]), .R(TRST_), .Q(
        DW4[22]) );
    zdffqrb DNT_DW4_Q_reg_21 ( .CK(DNT_DW4_n127), .D(ADI[21]), .R(TRST_), .Q(
        DW4[21]) );
    zdffqrb DNT_DW4_Q_reg_20 ( .CK(DNT_DW4_n127), .D(ADI[20]), .R(TRST_), .Q(
        DW4[20]) );
    zdffqrb DNT_DW4_Q_reg_19 ( .CK(DNT_DW4_n127), .D(ADI[19]), .R(TRST_), .Q(
        DW4[19]) );
    zdffqrb DNT_DW4_Q_reg_18 ( .CK(DNT_DW4_n127), .D(ADI[18]), .R(TRST_), .Q(
        DW4[18]) );
    zdffqrb DNT_DW4_Q_reg_17 ( .CK(DNT_DW4_n127), .D(ADI[17]), .R(TRST_), .Q(
        DW4[17]) );
    zdffqrb DNT_DW4_Q_reg_16 ( .CK(DNT_DW4_n127), .D(ADI[16]), .R(TRST_), .Q(
        DW4[16]) );
    zdffqrb DNT_DW4_Q_reg_15 ( .CK(DNT_DW4_n126), .D(ADI[15]), .R(TRST_), .Q(
        DW4[15]) );
    zdffqrb DNT_DW4_Q_reg_14 ( .CK(DNT_DW4_n126), .D(ADI[14]), .R(TRST_), .Q(
        DW4[14]) );
    zdffqrb DNT_DW4_Q_reg_13 ( .CK(DNT_DW4_n126), .D(ADI[13]), .R(TRST_), .Q(
        DW4[13]) );
    zdffqrb DNT_DW4_Q_reg_12 ( .CK(DNT_DW4_n126), .D(ADI[12]), .R(TRST_), .Q(
        DW4[12]) );
    zdffqrb DNT_DW4_Q_reg_11 ( .CK(DNT_DW4_n126), .D(ADI[11]), .R(TRST_), .Q(
        DW4[11]) );
    zdffqrb DNT_DW4_Q_reg_10 ( .CK(DNT_DW4_n126), .D(ADI[10]), .R(TRST_), .Q(
        DW4[10]) );
    zdffqrb DNT_DW4_Q_reg_9 ( .CK(DNT_DW4_n126), .D(ADI[9]), .R(TRST_), .Q(DW4
        [9]) );
    zdffqrb DNT_DW4_Q_reg_8 ( .CK(DNT_DW4_n126), .D(ADI[8]), .R(TRST_), .Q(DW4
        [8]) );
    zdffqrb DNT_DW4_Q_reg_7 ( .CK(DNT_DW4_n126), .D(ADI[7]), .R(TRST_), .Q(DW4
        [7]) );
    zdffqrb DNT_DW4_Q_reg_6 ( .CK(DNT_DW4_n126), .D(ADI[6]), .R(TRST_), .Q(DW4
        [6]) );
    zdffqrb DNT_DW4_Q_reg_5 ( .CK(DNT_DW4_n126), .D(ADI[5]), .R(TRST_), .Q(DW4
        [5]) );
    zdffqrb DNT_DW4_Q_reg_4 ( .CK(DNT_DW4_n126), .D(ADI[4]), .R(TRST_), .Q(DW4
        [4]) );
    zdffqrb DNT_DW4_Q_reg_3 ( .CK(DNT_DW4_n126), .D(ADI[3]), .R(TRST_), .Q(DW4
        [3]) );
    zdffqrb DNT_DW4_Q_reg_2 ( .CK(DNT_DW4_n126), .D(ADI[2]), .R(TRST_), .Q(DW4
        [2]) );
    zdffqrb DNT_DW4_Q_reg_1 ( .CK(DNT_DW4_n126), .D(ADI[1]), .R(TRST_), .Q(DW4
        [1]) );
    zdffqrb DNT_DW4_Q_reg_0 ( .CK(DNT_DW4_n126), .D(ADI[0]), .R(TRST_), .Q(DW4
        [0]) );
    zbfb DNT_DW4_U80 ( .A(FLOPS_CLK_8), .Y(DNT_DW4_n126) );
    zbfb DNT_DW4_U81 ( .A(FLOPS_CLK_8), .Y(DNT_DW4_n127) );
endmodule


module HS_FMTIMER ( CLK60M, TRST_, FLADJ, REDUCE, EOF1, EOF2, PRESOF, FRNUM, 
    PCICLK, MAXLEN, SOFV, ADI, WR_FRNUM, RUN, HCHALT, FRLSTSIZE, SOFGEN, 
    EHCISLEEP, EHCIRESTART, START_EVENT, FROZEN, ROLLOVER_S, INTTHRESHOLD, 
    ITDIOCINT1, ITDIOCINT2, SITDIOCINT1, SITDIOCINT2, USBINT, ERRINT, INTASYNC, 
    QHIOCINT1, QHIOCINT2, QHIOCINT3, QHIOCINT4, QHERRINT1, QHERRINT2, 
    QHERRINT3, QHERRINT4, QHASYNCINT, ASYNCINT, GEN_PERR, ASYNC_ACT, SWDBG, 
    MAC_EOT, EHCI_MAC_EOT, EHCI_DBG_MAC_EOT, HSERR_S, FRNUM_PCLK, FRNUM_AD, 
    PRESOF_EVAL, HCI_PRESOF, LTINT_PCLK, FRNUM_PCLK_LATCH, CMDSTART, TXSOF, 
    SLEEPTIME_SEL, ATPG_ENI );
input  [5:0] FLADJ;
output [13:0] FRNUM;
input  [1:0] FRLSTSIZE;
output [13:0] FRNUM_PCLK;
input  [10:0] MAXLEN;
output [10:0] SOFV;
input  [31:0] ADI;
input  [7:0] INTTHRESHOLD;
output [13:0] FRNUM_AD;
input  CLK60M, TRST_, REDUCE, PCICLK, WR_FRNUM, RUN, HCHALT, EHCISLEEP, 
    START_EVENT, FROZEN, ITDIOCINT1, ITDIOCINT2, SITDIOCINT1, SITDIOCINT2, 
    USBINT, ERRINT, INTASYNC, QHIOCINT1, QHIOCINT2, QHIOCINT3, QHIOCINT4, 
    QHERRINT1, QHERRINT2, QHERRINT3, QHERRINT4, QHASYNCINT, GEN_PERR, 
    ASYNC_ACT, SWDBG, MAC_EOT, EHCI_DBG_MAC_EOT, HSERR_S, PRESOF_EVAL, 
    HCI_PRESOF, CMDSTART, TXSOF, SLEEPTIME_SEL, ATPG_ENI;
output EOF1, EOF2, PRESOF, SOFGEN, EHCIRESTART, ROLLOVER_S, ASYNCINT, 
    EHCI_MAC_EOT, LTINT_PCLK, FRNUM_PCLK_LATCH;
    wire CMDTXSOF, FRNUM730_13, SOFV769_3, TMCNT_EN1460, TMCNT1530_2, SPAREO6, 
        FRNUM730_7, TMCNT1516_10, TMCNT_12, FRNUM_PCLK575_9, n1131_31, 
        FRNUMNXT_T_9, FMREMN_5, TMCNT1516_5, EOF11263, SOFGEN1084, 
        FMREMN1078_8, FMREMNXT957_7, FRNUMNXT_T_11, val313_4, ROLLOVER_S_T633, 
        FMINTV_3, TMCNT_2, LTINT_CK, PRESOF_CAL_6, n1131_23, FRNUM_W484_13, 
        FMREMNXT_4, FRNUM_PCLK575_0, EHCIRESTART1600, FRNUM_W484_7, 
        FRAMECHG_2T, b1610_1, FRNUM_W_2, FMREMN1078_1, FRNUMNXT_T_7, EOF21267, 
        FMREMN1078_6, FRNUM_W_5, FMREMNXT957_9, SPAREO0_, FRNUM_W484_0, 
        FRNUM_PCLK575_7, n1131_24, PRESOF_CAL_1, FMREMNXT_3, SPAREO8, 
        FRNUM730_9, FRNUM_W_10, TMCNT_EN, TMCNT_5, FMINTV_4, FRCHGCHKBIT_T, 
        FRNUM_PCLK575_13, FMREMN_2, TMCNT1516_2, START_EVENT_3T, FMREMN_11, 
        FRNUM_W484_9, TMCNT1530_5, PRESOF_CAL_8, SOFV769_4, FRNUM730_0, 
        SPAREO1, FRNUM_W_11, FMINTV_5, TMCNT_4, FRNUM_PCLK575_12, n1131_25, 
        FRCHGCHKBIT, FMREMNXT_2, SPAREO9, FRNUM730_8, WR_FRNUMT, WR_FRNUMT_2T, 
        FRNUM_W484_1, FRNUM_PCLK575_6, FRNUMNXT_T_6, FRAMECHG1090, 
        FMREMN1078_7, FRNUM_W_4, FMREMNXT957_12, FMREMNXT957_8, PRESOF1203, 
        PRESOF_CAL_9, TMCNT1530_4, SOFV769_10, SOFV769_5, EHCI_MAC_EOT_PCLK, 
        FRNUM730_1, SPAREO0, HSERR_S_T, FMREMN1078_12, FMREMN_10, FRNUM_W484_8, 
        FMREMN_3, TMCNT1516_3, FMREMNXT957_1, FRNUMNXT_T_8, FMREMN_4, 
        TMCNT1516_4, EOF11262, FMREMN1078_9, FMREMNXT957_6, FRNUM_PCLK575_8, 
        n1131_30, SOFV769_2, TMCNT1530_12, TMCNT1530_3, SPAREO7, TMCNT1516_11, 
        FRNUM730_6, FROZSYNC, n1311, FRNUM_W_3, FRNUM730_12, FRNUMNXT_T_1, 
        LTINT, FMREMN1078_0, CMDTXSOF_3T, FRNUM_PCLK575_1, FRNUM_W484_6, 
        RSTREMAIN_, PRESOF_CAL_7, CMDTXSOF1868, FRNUM_W484_12, FMREMNXT_5, 
        FRNUMNXT_T_10, LTINT_PCLK1831, START_EVENT_T, ROLLCHKBIT, FMREMNXT_12, 
        FMINTV_2, TMCNT_3, TMCNT_8, FRNUM730_10, FRNUM730_4, CMDTXSOF_2T, 
        SPAREO5, TMCNT1530_10, TMCNT1530_1, SOFV769_0, n1131_29, TMCNT_11, 
        START_EVENT_SYNC1423, FRNUM_W_8, FMREMNXT957_4, FMREMN_6, TMCNT1516_6, 
        TMCNT_1, PRESOF_CAL_10, FMREMNXT_10, FRAMECHG, FRNUMNXT_T_12, 
        FMREMNXT_7, START_EVENT_SYNC, FRNUM_W484_10, SOFV769_9, TMCNT1530_8, 
        PRESOF_CAL_5, FRNUM_W484_4, FRNUM_PCLK575_3, FMREMN1078_2, FRNUM_W_6, 
        FRNUM_W_1, FRNUMNXT_T_3, FMREMNXT957_10, FMREMN1078_5, FRNUMNXT_T_4, 
        FMREMN_8, TMCNT1516_8, FRNUM_PCLK575_4, FRNUM_W484_3, ROLLCHKBIT_T, 
        FMREMNXT_0, FRNUM_W_13, PRESOF_CAL_2, n1131_27, FRNUM_PCLK575_10, 
        TMCNT_6, FMINTV_7, FMREMNXT957_3, FMREMN_1, TMCNT1516_1, FMREMN_12, 
        FMREMN1078_10, SPAREO2, FMREMNXT_9, FRAMECHG_T, FRNUM730_3, SOFV769_7, 
        WR_FRNUMT_3T, TMCNT1530_6, FRNUM_W_12, FRNUM_PCLK575_11, PRESOF1187, 
        FMINTV_6, TMCNT_7, FMREMNXT_1, START_EVENT_2T, c1612_1, PRESOF_CAL_3, 
        n1131_26, FRNUM_PCLK575_5, FRNUM_W484_2, FMREMNXT957_11, FRNUM_W_7, 
        FMREMN1078_4, FRNUMNXT_T_5, FMREMN_9, TMCNT1516_9, SPAREO3, FMREMNXT_8, 
        FRNUM730_2, SPAREO1_, SOFV769_6, TMCNT1530_7, FRCHGCHKBIT_2T, 
        WR_FRNUMT_T, FMREMN1078_11, FRNUM_W_9, FMREMNXT957_2, TMCNT1516_0, 
        HSERR_S_2T, n1309, FMREMNXT957_5, FMREMN_7, TMCNT1516_7, WR_FRNUMT393, 
        TMCNT_10, TMCNT1516_12, FRNUM730_5, SPAREO4, TMCNT1530_11, TMCNT1530_0, 
        SOFV769_1, n1131_28, TMCNT_9, FRNUM730_11, FMREMN1078_3, FRNUM_W_0, 
        FRNUMNXT_T_2, ROLLOVER_S_T, FRNUM_W484_5, FRNUM_PCLK575_2, FMREMNXT_6, 
        FRNUM_W484_11, SOFV769_8, PRESOF_CAL_4, TMCNT1530_9, CMDTXSOF_T, 
        FMINTV_1, TMCNT_0, PRESOF_CAL_11, FMREMNXT_11, FRNUMNXT_T_13, n2325, 
        n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, 
        add_60_carry_6, add_60_carry_2, add_60_carry_5, add_60_carry_4, 
        add_60_carry_3, add_175_carry_8, add_175_carry_12, add_175_carry_6, 
        add_175_carry_13, add_175_carry_7, add_175_carry_9, add_175_carry_2, 
        add_175_carry_11, add_175_carry_5, add_175_carry_10, add_175_carry_4, 
        add_175_carry_3, sub_325_carry_12, sub_325_carry_8, sub_325_carry_1, 
        sub_325_carry_7, sub_325_carry_6, sub_325_carry_11, sub_325_carry_9, 
        sub_325_carry_2, sub_325_carry_10, sub_325_carry_5, sub_325_carry_4, 
        sub_325_carry_3, add_378_carry_8, add_378_carry_1, add_378_carry_7, 
        add_378_carry_6, add_378_carry_9, add_378_carry_2, add_378_carry_10, 
        add_378_carry_5, add_378_carry_4, add_378_carry_3, add_378_2_carry_8, 
        add_378_2_carry_7, add_378_2_carry_6, add_378_2_carry_5, 
        add_378_2_carry_4, add_378_2_carry_3, n2346, n2347, n2348, n2349, 
        n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, 
        n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
        n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, 
        n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, 
        n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, 
        n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, 
        n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, 
        n2420, n2421, n2422, n2423, n2424, n2425, add_500_carry_8, 
        add_500_carry_12, add_500_carry_6, add_500_carry_7, add_500_carry_9, 
        add_500_carry_2, add_500_carry_11, add_500_carry_5, add_500_carry_10, 
        add_500_carry_4, add_500_carry_3, n2426, n2427, n2428, n2429, n2430, 
        n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, 
        n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
        n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
        n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, 
        n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, 
        n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
        n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
        n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, 
        n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
        n2521, n2523, n2524, n2525;
    assign FRNUM_AD[13] = 1'b0;
    zaoi211b SPARE542 ( .A(SPAREO0), .B(WR_FRNUMT_2T), .C(SPAREO1_), .D(1'b0), 
        .Y(SPAREO2) );
    zoai21b SPARE545 ( .A(SPAREO1), .B(RSTREMAIN_), .C(SPAREO9), .Y(SPAREO3)
         );
    zoai21b SPARE544 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zmux21hb DNTCK ( .A(LTINT), .B(CLK60M), .S(ATPG_ENI), .Y(LTINT_CK) );
    zaoi211b SPARE543 ( .A(SPAREO4), .B(FRCHGCHKBIT), .C(SPAREO6), .D(1'b0), 
        .Y(SPAREO8) );
    zivb SPARE548 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE541 ( .CK(CLK60M), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    znr3b SPARE546 ( .A(SPAREO2), .B(LTINT), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE547 ( .A(SPAREO4), .Y(SPAREO5) );
    znd3b SPARE549 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE540 ( .CK(CLK60M), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd2b U742 ( .A(FMREMNXT_1), .B(n2372), .Y(n2365) );
    znd2b U743 ( .A(FMREMNXT_0), .B(n2332), .Y(n2363) );
    zivb U744 ( .A(PRESOF_CAL_1), .Y(n2372) );
    znd2b U745 ( .A(FMREMNXT_3), .B(n2370), .Y(n2358) );
    znd2b U746 ( .A(FMREMNXT_2), .B(n2373), .Y(n2364) );
    znd3b U747 ( .A(n2360), .B(n2362), .C(n2361), .Y(n2359) );
    znd2b U748 ( .A(PRESOF_CAL_1), .B(n2374), .Y(n2360) );
    znd2b U749 ( .A(n2363), .B(n2365), .Y(n2362) );
    znd2b U750 ( .A(PRESOF_CAL_2), .B(n2412), .Y(n2361) );
    zivb U751 ( .A(PRESOF_CAL_3), .Y(n2370) );
    zivb U752 ( .A(PRESOF_CAL_2), .Y(n2373) );
    znd2b U753 ( .A(FMREMNXT_5), .B(n2368), .Y(n2352) );
    znd2b U754 ( .A(FMREMNXT_4), .B(n2371), .Y(n2357) );
    znd3b U755 ( .A(n2354), .B(n2356), .C(n2355), .Y(n2353) );
    znd2b U756 ( .A(PRESOF_CAL_3), .B(n2396), .Y(n2354) );
    znd3b U757 ( .A(n2359), .B(n2364), .C(n2358), .Y(n2356) );
    znd2b U758 ( .A(PRESOF_CAL_4), .B(n2419), .Y(n2355) );
    zivb U759 ( .A(PRESOF_CAL_5), .Y(n2368) );
    zivb U760 ( .A(PRESOF_CAL_4), .Y(n2371) );
    znd2b U761 ( .A(FMREMNXT_7), .B(n2387), .Y(n2346) );
    znd2b U762 ( .A(FMREMNXT_6), .B(n2369), .Y(n2351) );
    zivb U763 ( .A(PRESOF_CAL_6), .Y(n2369) );
    znd3b U764 ( .A(n2348), .B(n2350), .C(n2349), .Y(n2347) );
    znd2b U765 ( .A(PRESOF_CAL_5), .B(n2399), .Y(n2348) );
    znd3b U766 ( .A(n2353), .B(n2357), .C(n2352), .Y(n2350) );
    znd2b U767 ( .A(PRESOF_CAL_6), .B(n2424), .Y(n2349) );
    znr2b U768 ( .A(FMREMNXT_8), .B(n2389), .Y(n2390) );
    znr2b U769 ( .A(FMREMNXT_7), .B(n2387), .Y(n2388) );
    zivb U770 ( .A(PRESOF_CAL_8), .Y(n2389) );
    zivb U771 ( .A(PRESOF_CAL_7), .Y(n2387) );
    znr2b U772 ( .A(FMREMNXT_9), .B(n2384), .Y(n2385) );
    znr2b U773 ( .A(FMREMNXT_10), .B(n2382), .Y(n2383) );
    znd2b U774 ( .A(FMREMNXT_9), .B(n2384), .Y(n2379) );
    zaoi21b U775 ( .A(n2367), .B(n2366), .C(n2392), .Y(n2380) );
    znr2b U776 ( .A(n2388), .B(n2390), .Y(n2367) );
    znd3b U777 ( .A(n2347), .B(n2351), .C(n2346), .Y(n2366) );
    znr2b U778 ( .A(PRESOF_CAL_8), .B(n2391), .Y(n2392) );
    zivb U779 ( .A(PRESOF_CAL_10), .Y(n2382) );
    zivb U780 ( .A(PRESOF_CAL_9), .Y(n2384) );
    znr2b U781 ( .A(n2430), .B(n2434), .Y(n2431) );
    znd2b U782 ( .A(TMCNT_4), .B(TMCNT_5), .Y(n2430) );
    znd2b U783 ( .A(n2432), .B(n2433), .Y(n2428) );
    znr2b U784 ( .A(TMCNT_0), .B(TMCNT_2), .Y(n2432) );
    znr2b U785 ( .A(TMCNT_3), .B(TMCNT_1), .Y(n2433) );
    znr2b U786 ( .A(FMREMNXT_11), .B(n2375), .Y(n2376) );
    zivb U787 ( .A(PRESOF_CAL_11), .Y(n2375) );
    znr3b U788 ( .A(n2378), .B(n2386), .C(n2381), .Y(n2377) );
    znr2b U789 ( .A(PRESOF_CAL_11), .B(n2403), .Y(n2378) );
    znr2b U790 ( .A(PRESOF_CAL_10), .B(n2410), .Y(n2386) );
    zaoi211b U791 ( .A(n2380), .B(n2379), .C(n2383), .D(n2385), .Y(n2381) );
    znd3b U792 ( .A(n2397), .B(n2396), .C(n2419), .Y(n2398) );
    znd3b U793 ( .A(FMREMNXT_0), .B(FMREMNXT_1), .C(FMREMNXT_2), .Y(n2397) );
    zxo2b U794 ( .A(FRNUM[1]), .B(FRNUMNXT_T_1), .Y(n2490) );
    znd2b U795 ( .A(n2429), .B(n2427), .Y(n2426) );
    znr2b U796 ( .A(TMCNT_7), .B(TMCNT_8), .Y(n2429) );
    znd2b U797 ( .A(n2428), .B(n2431), .Y(n2427) );
    znd2b U798 ( .A(n2410), .B(n2409), .Y(n2411) );
    znd2b U799 ( .A(n2404), .B(n2403), .Y(n2405) );
    zaoi21b U800 ( .A(n2413), .B(n2412), .C(n2396), .Y(n2414) );
    znr2b U801 ( .A(FMREMNXT_1), .B(FMREMNXT_0), .Y(n2413) );
    zaoi21b U802 ( .A(FMREMNXT_1), .B(FMREMNXT_0), .C(FMREMNXT_2), .Y(n2417)
         );
    znr2b U803 ( .A(FMREMNXT_11), .B(FMREMNXT_12), .Y(n2418) );
    znr2b U804 ( .A(FMREMNXT_10), .B(FMREMNXT_3), .Y(n2422) );
    znr2b U805 ( .A(FMREMNXT_9), .B(FMREMNXT_8), .Y(n2420) );
    zxn2b sub_325_U1_A_12 ( .A(FMREMN_12), .B(sub_325_carry_12), .Y(
        FMREMNXT957_12) );
    zor2b sub_325_U1_B_11 ( .A(FMREMN_11), .B(sub_325_carry_11), .Y(
        sub_325_carry_12) );
    zxn2b sub_325_U1_A_6 ( .A(FMREMN_6), .B(sub_325_carry_6), .Y(FMREMNXT957_6
        ) );
    zor2b sub_325_U1_B_5 ( .A(FMREMN_5), .B(sub_325_carry_5), .Y(
        sub_325_carry_6) );
    zxn2b sub_325_U1_A_1 ( .A(FMREMN_1), .B(sub_325_carry_1), .Y(FMREMNXT957_1
        ) );
    znr2b U806 ( .A(n2393), .B(FMREMNXT_12), .Y(PRESOF1187) );
    znr2b U807 ( .A(HCI_PRESOF), .B(n2505), .Y(n2518) );
    zxn2b sub_325_U1_A_8 ( .A(FMREMN_8), .B(sub_325_carry_8), .Y(FMREMNXT957_8
        ) );
    zor2b sub_325_U1_B_7 ( .A(FMREMN_7), .B(sub_325_carry_7), .Y(
        sub_325_carry_8) );
    zxn2b sub_325_U1_A_9 ( .A(FMREMN_9), .B(sub_325_carry_9), .Y(FMREMNXT957_9
        ) );
    zor2b sub_325_U1_B_8 ( .A(FMREMN_8), .B(sub_325_carry_8), .Y(
        sub_325_carry_9) );
    znd3b U808 ( .A(n2409), .B(n2395), .C(n2394), .Y(n2401) );
    znr2b U809 ( .A(FMREMNXT_10), .B(FMREMNXT_8), .Y(n2395) );
    znr2b U810 ( .A(FMREMNXT_11), .B(FMREMNXT_12), .Y(n2394) );
    znr2b U811 ( .A(n2400), .B(n2406), .Y(n2402) );
    zxo2b U812 ( .A(n2511), .B(n2474), .Y(n2480) );
    zan2b U813 ( .A(n2475), .B(n2476), .Y(n2474) );
    zoa22b U814 ( .A(n2475), .B(n2476), .C(n2487), .D(n2512), .Y(n2479) );
    zivb U815 ( .A(INTTHRESHOLD[2]), .Y(n2512) );
    zor2b U816 ( .A(n2521), .B(n2513), .Y(n2478) );
    zan3b U817 ( .A(n2485), .B(n2520), .C(n2491), .Y(n2477) );
    zivb U818 ( .A(INTTHRESHOLD[7]), .Y(n2520) );
    zivb U819 ( .A(INTTHRESHOLD[5]), .Y(n2513) );
    zxo2b U820 ( .A(n2495), .B(FRNUM[5]), .Y(n2494) );
    zmux21lb U821 ( .A(INTTHRESHOLD[0]), .B(n2489), .S(INTTHRESHOLD[1]), .Y(
        n2481) );
    zan2b U822 ( .A(n2490), .B(n2491), .Y(n2489) );
    zivb U823 ( .A(INTTHRESHOLD[0]), .Y(n2491) );
    zxo2b U824 ( .A(n2493), .B(FRNUM[6]), .Y(n2492) );
    zor2b U825 ( .A(INTTHRESHOLD[2]), .B(n2508), .Y(n2509) );
    zivb U826 ( .A(n2509), .Y(n2521) );
    zor2b U827 ( .A(INTTHRESHOLD[0]), .B(INTTHRESHOLD[1]), .Y(n2510) );
    zivb U828 ( .A(n2510), .Y(n2476) );
    zan2b U829 ( .A(n2487), .B(n2488), .Y(n2486) );
    zivb U830 ( .A(n2508), .Y(n2487) );
    zor2b U831 ( .A(INTTHRESHOLD[3]), .B(INTTHRESHOLD[4]), .Y(n2508) );
    zxo2b U832 ( .A(FRNUM[2]), .B(FRNUMNXT_T_2), .Y(n2488) );
    zan3b U833 ( .A(n2484), .B(INTTHRESHOLD[4]), .C(n2485), .Y(n2483) );
    zxo2b U834 ( .A(FRNUM[4]), .B(FRNUMNXT_T_4), .Y(n2484) );
    zivb U835 ( .A(INTTHRESHOLD[3]), .Y(n2485) );
    zxn2b sub_325_U1_A_7 ( .A(FMREMN_7), .B(sub_325_carry_7), .Y(FMREMNXT957_7
        ) );
    zor2b sub_325_U1_B_6 ( .A(FMREMN_6), .B(sub_325_carry_6), .Y(
        sub_325_carry_7) );
    zxn2b sub_325_U1_A_11 ( .A(FMREMN_11), .B(sub_325_carry_11), .Y(
        FMREMNXT957_11) );
    zor2b sub_325_U1_B_10 ( .A(FMREMN_10), .B(sub_325_carry_10), .Y(
        sub_325_carry_11) );
    zxn2b sub_325_U1_A_5 ( .A(FMREMN_5), .B(sub_325_carry_5), .Y(FMREMNXT957_5
        ) );
    zor2b sub_325_U1_B_4 ( .A(FMREMN_4), .B(sub_325_carry_4), .Y(
        sub_325_carry_5) );
    zxn2b sub_325_U1_A_2 ( .A(FMREMN_2), .B(sub_325_carry_2), .Y(FMREMNXT957_2
        ) );
    zor2b sub_325_U1_B_1 ( .A(FMREMN_1), .B(sub_325_carry_1), .Y(
        sub_325_carry_2) );
    zan2b U836 ( .A(FRNUM[11]), .B(n2504), .Y(n2516) );
    zan2b U837 ( .A(FRLSTSIZE[0]), .B(FRNUM[12]), .Y(n2517) );
    znd2b U838 ( .A(n2436), .B(n2435), .Y(b1610_1) );
    znr3b U839 ( .A(TMCNT_12), .B(TMCNT_10), .C(TMCNT_11), .Y(n2436) );
    znd2b U840 ( .A(TMCNT_9), .B(n2426), .Y(n2435) );
    znd3b U841 ( .A(n2439), .B(n2438), .C(n2437), .Y(c1612_1) );
    znr2b U842 ( .A(TMCNT_9), .B(TMCNT_8), .Y(n2439) );
    znr2b U843 ( .A(TMCNT_7), .B(TMCNT_10), .Y(n2438) );
    znr3b U844 ( .A(TMCNT_6), .B(TMCNT_11), .C(TMCNT_12), .Y(n2437) );
    zxn2b sub_325_U1_A_3 ( .A(FMREMN_3), .B(sub_325_carry_3), .Y(FMREMNXT957_3
        ) );
    zor2b sub_325_U1_B_2 ( .A(FMREMN_2), .B(sub_325_carry_2), .Y(
        sub_325_carry_3) );
    znd3b U845 ( .A(n2407), .B(n2408), .C(n2406), .Y(n2415) );
    znr3b U846 ( .A(FMREMNXT_5), .B(n2414), .C(n2405), .Y(n2407) );
    znr3b U847 ( .A(FMREMNXT_4), .B(n2411), .C(FMREMNXT_8), .Y(n2408) );
    znr2b U848 ( .A(n2421), .B(n2416), .Y(n2425) );
    znd3b U849 ( .A(n2420), .B(n2422), .C(n2419), .Y(n2421) );
    znd3b U850 ( .A(n2418), .B(n2417), .C(n2399), .Y(n2416) );
    zxn2b sub_325_U1_A_10 ( .A(FMREMN_10), .B(sub_325_carry_10), .Y(
        FMREMNXT957_10) );
    zor2b sub_325_U1_B_9 ( .A(FMREMN_9), .B(sub_325_carry_9), .Y(
        sub_325_carry_10) );
    znr2b U851 ( .A(FROZSYNC), .B(n2515), .Y(n2325) );
    zivb U852 ( .A(n2515), .Y(n2514) );
    zxn2b sub_325_U1_A_4 ( .A(FMREMN_4), .B(sub_325_carry_4), .Y(FMREMNXT957_4
        ) );
    zor2b sub_325_U1_B_3 ( .A(FMREMN_3), .B(sub_325_carry_3), .Y(
        sub_325_carry_4) );
    zan2b U853 ( .A(n2472), .B(n2473), .Y(n2471) );
    zan2b U854 ( .A(RSTREMAIN_), .B(FMREMNXT_0), .Y(FMREMN1078_0) );
    zmux21hb U855 ( .A(FRNUM[0]), .B(FRNUM_AD[0]), .S(n2519), .Y(
        FRNUM_PCLK575_0) );
    zmux21hb U856 ( .A(FRNUM[1]), .B(FRNUM_AD[1]), .S(n2519), .Y(
        FRNUM_PCLK575_1) );
    zmux21hb U857 ( .A(FRNUM[2]), .B(FRNUM_AD[2]), .S(n2519), .Y(
        FRNUM_PCLK575_2) );
    zmux21hb U858 ( .A(FRNUM[3]), .B(FRNUM_AD[3]), .S(n2519), .Y(
        FRNUM_PCLK575_3) );
    zmux21hb U859 ( .A(FRNUM[4]), .B(FRNUM_AD[4]), .S(n2519), .Y(
        FRNUM_PCLK575_4) );
    zmux21hb U860 ( .A(FRNUM[5]), .B(FRNUM_AD[5]), .S(n2519), .Y(
        FRNUM_PCLK575_5) );
    zmux21hb U861 ( .A(FRNUM[6]), .B(FRNUM_AD[6]), .S(n2519), .Y(
        FRNUM_PCLK575_6) );
    zmux21hb U862 ( .A(FRNUM[7]), .B(FRNUM_AD[7]), .S(n2519), .Y(
        FRNUM_PCLK575_7) );
    zmux21hb U863 ( .A(FRNUM[8]), .B(FRNUM_AD[8]), .S(n2519), .Y(
        FRNUM_PCLK575_8) );
    zmux21hb U864 ( .A(FRNUM[9]), .B(FRNUM_AD[9]), .S(n2519), .Y(
        FRNUM_PCLK575_9) );
    zmux21hb U865 ( .A(FRNUM[10]), .B(FRNUM_AD[10]), .S(n2519), .Y(
        FRNUM_PCLK575_10) );
    zan2b U866 ( .A(FRNUM_W_13), .B(n2453), .Y(FRNUM_W484_13) );
    zmux21hb U867 ( .A(FRNUM_W_12), .B(ADI[12]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_12) );
    zmux21hb U868 ( .A(FRNUM_W_11), .B(ADI[11]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_11) );
    zmux21hb U869 ( .A(FRNUM_W_10), .B(ADI[10]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_10) );
    zmux21hb U870 ( .A(FRNUM_W_9), .B(ADI[9]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_9) );
    zmux21hb U871 ( .A(FRNUM_W_8), .B(ADI[8]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_8) );
    zmux21hb U872 ( .A(FRNUM_W_7), .B(ADI[7]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_7) );
    zmux21hb U873 ( .A(FRNUM_W_6), .B(ADI[6]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_6) );
    zmux21hb U874 ( .A(FRNUM_W_5), .B(ADI[5]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_5) );
    zmux21hb U875 ( .A(FRNUM_W_4), .B(ADI[4]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_4) );
    zmux21hb U876 ( .A(FRNUM_W_3), .B(ADI[3]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_3) );
    zmux21hb U877 ( .A(FRNUM_W_2), .B(ADI[2]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_2) );
    zmux21hb U878 ( .A(FRNUM_W_1), .B(ADI[1]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_1) );
    zmux21hb U879 ( .A(FRNUM_W_0), .B(ADI[0]), .S(WR_FRNUMT393), .Y(
        FRNUM_W484_0) );
    zmux21hb U880 ( .A(FRNUM[13]), .B(FRNUM_PCLK[13]), .S(n2519), .Y(
        FRNUM_PCLK575_13) );
    zmux21lb U881 ( .A(n2499), .B(n2506), .S(n2519), .Y(FRNUM_PCLK575_12) );
    zmux21lb U882 ( .A(n2500), .B(n2507), .S(n2519), .Y(FRNUM_PCLK575_11) );
    zxo2b U883 ( .A(add_175_carry_13), .B(FRNUM[13]), .Y(FRNUMNXT_T_13) );
    zhadrb add_175_U1_1_12 ( .A(FRNUM[12]), .B(add_175_carry_12), .CO(
        add_175_carry_13), .S(FRNUMNXT_T_12) );
    zhadrb add_175_U1_1_11 ( .A(FRNUM[11]), .B(add_175_carry_11), .CO(
        add_175_carry_12), .S(FRNUMNXT_T_11) );
    zhadrb add_175_U1_1_10 ( .A(FRNUM[10]), .B(add_175_carry_10), .CO(
        add_175_carry_11), .S(FRNUMNXT_T_10) );
    zhadrb add_175_U1_1_9 ( .A(FRNUM[9]), .B(add_175_carry_9), .CO(
        add_175_carry_10), .S(FRNUMNXT_T_9) );
    zhadrb add_175_U1_1_8 ( .A(FRNUM[8]), .B(add_175_carry_8), .CO(
        add_175_carry_9), .S(FRNUMNXT_T_8) );
    zhadrb add_175_U1_1_7 ( .A(FRNUM[7]), .B(add_175_carry_7), .CO(
        add_175_carry_8), .S(FRNUMNXT_T_7) );
    zhadrb add_175_U1_1_6 ( .A(FRNUM[6]), .B(add_175_carry_6), .CO(
        add_175_carry_7), .S(FRNUMNXT_T_6) );
    zivb U884 ( .A(FRNUMNXT_T_6), .Y(n2493) );
    zhadrb add_175_U1_1_5 ( .A(FRNUM[5]), .B(add_175_carry_5), .CO(
        add_175_carry_6), .S(FRNUMNXT_T_5) );
    zivb U885 ( .A(FRNUMNXT_T_5), .Y(n2495) );
    zhadrb add_175_U1_1_4 ( .A(FRNUM[4]), .B(add_175_carry_4), .CO(
        add_175_carry_5), .S(FRNUMNXT_T_4) );
    zhadrb add_175_U1_1_3 ( .A(FRNUM[3]), .B(add_175_carry_3), .CO(
        add_175_carry_4), .S(FRNUMNXT_T_3) );
    zhadrb add_175_U1_1_2 ( .A(FRNUM[2]), .B(add_175_carry_2), .CO(
        add_175_carry_3), .S(FRNUMNXT_T_2) );
    zhadrb add_175_U1_1_1 ( .A(FRNUM[1]), .B(FRNUM[0]), .CO(add_175_carry_2), 
        .S(FRNUMNXT_T_1) );
    zmux21hb U886 ( .A(FRNUM[13]), .B(SOFV[10]), .S(n2330), .Y(SOFV769_10) );
    zmux21hb U887 ( .A(FRNUM[12]), .B(SOFV[9]), .S(n2330), .Y(SOFV769_9) );
    zmux21hb U888 ( .A(FRNUM[11]), .B(SOFV[8]), .S(n2330), .Y(SOFV769_8) );
    zmux21hb U889 ( .A(FRNUM[10]), .B(SOFV[7]), .S(n2330), .Y(SOFV769_7) );
    zmux21hb U890 ( .A(FRNUM[9]), .B(SOFV[6]), .S(n2330), .Y(SOFV769_6) );
    zmux21hb U891 ( .A(FRNUM[8]), .B(SOFV[5]), .S(n2330), .Y(SOFV769_5) );
    zmux21hb U892 ( .A(FRNUM[7]), .B(SOFV[4]), .S(n2330), .Y(SOFV769_4) );
    zmux21hb U893 ( .A(FRNUM[6]), .B(SOFV[3]), .S(n2330), .Y(SOFV769_3) );
    zmux21hb U894 ( .A(FRNUM[5]), .B(SOFV[2]), .S(n2330), .Y(SOFV769_2) );
    zmux21hb U895 ( .A(FRNUM[4]), .B(SOFV[1]), .S(n2330), .Y(SOFV769_1) );
    zmux21hb U896 ( .A(FRNUM[3]), .B(SOFV[0]), .S(n2330), .Y(SOFV769_0) );
    zxo2b U897 ( .A(add_500_carry_12), .B(TMCNT_12), .Y(TMCNT1516_12) );
    zhadrb add_500_U1_1_11 ( .A(TMCNT_11), .B(add_500_carry_11), .CO(
        add_500_carry_12), .S(TMCNT1516_11) );
    zhadrb add_500_U1_1_10 ( .A(TMCNT_10), .B(add_500_carry_10), .CO(
        add_500_carry_11), .S(TMCNT1516_10) );
    zhadrb add_500_U1_1_9 ( .A(TMCNT_9), .B(add_500_carry_9), .CO(
        add_500_carry_10), .S(TMCNT1516_9) );
    zhadrb add_500_U1_1_8 ( .A(TMCNT_8), .B(add_500_carry_8), .CO(
        add_500_carry_9), .S(TMCNT1516_8) );
    zhadrb add_500_U1_1_7 ( .A(TMCNT_7), .B(add_500_carry_7), .CO(
        add_500_carry_8), .S(TMCNT1516_7) );
    zhadrb add_500_U1_1_6 ( .A(TMCNT_6), .B(add_500_carry_6), .CO(
        add_500_carry_7), .S(TMCNT1516_6) );
    zhadrb add_500_U1_1_5 ( .A(TMCNT_5), .B(add_500_carry_5), .CO(
        add_500_carry_6), .S(TMCNT1516_5) );
    zhadrb add_500_U1_1_4 ( .A(TMCNT_4), .B(add_500_carry_4), .CO(
        add_500_carry_5), .S(TMCNT1516_4) );
    zhadrb add_500_U1_1_3 ( .A(TMCNT_3), .B(add_500_carry_3), .CO(
        add_500_carry_4), .S(TMCNT1516_3) );
    zhadrb add_500_U1_1_2 ( .A(TMCNT_2), .B(add_500_carry_2), .CO(
        add_500_carry_3), .S(TMCNT1516_2) );
    zhadrb add_500_U1_1_1 ( .A(TMCNT_1), .B(TMCNT_0), .CO(add_500_carry_2), 
        .S(TMCNT1516_1) );
    zan2b U898 ( .A(RSTREMAIN_), .B(FMREMNXT_12), .Y(FMREMN1078_12) );
    zivb U899 ( .A(FMREMNXT_12), .Y(n2404) );
    zan2b U900 ( .A(RSTREMAIN_), .B(FMREMNXT_6), .Y(FMREMN1078_6) );
    zxo2b U901 ( .A(ROLLCHKBIT), .B(ROLLCHKBIT_T), .Y(ROLLOVER_S_T633) );
    zor2b U902 ( .A(FMREMNXT_1), .B(n2450), .Y(FMREMN1078_1) );
    zivb U903 ( .A(FMREMNXT_1), .Y(n2374) );
    zivb U904 ( .A(n2453), .Y(WR_FRNUMT393) );
    znd3b U905 ( .A(HCHALT), .B(WR_FRNUM), .C(n2473), .Y(n2453) );
    zivb U906 ( .A(RUN), .Y(n2473) );
    znd2b U907 ( .A(n2454), .B(RSTREMAIN_), .Y(PRESOF1203) );
    zmux21lb U908 ( .A(n2518), .B(PRESOF1187), .S(PRESOF_EVAL), .Y(n2454) );
    zan2b U909 ( .A(RSTREMAIN_), .B(FMREMNXT_8), .Y(FMREMN1078_8) );
    zivb U910 ( .A(FMREMNXT_8), .Y(n2391) );
    zcx4b U911 ( .A(TMCNT_EN), .B(EHCISLEEP), .C(START_EVENT_SYNC), .D(n2452), 
        .Y(TMCNT_EN1460) );
    zor2b U912 ( .A(EHCIRESTART), .B(PRESOF), .Y(n2452) );
    zan2b U913 ( .A(RSTREMAIN_), .B(FMREMNXT_9), .Y(FMREMN1078_9) );
    zor2b U914 ( .A(EOF11263), .B(n2450), .Y(EOF11262) );
    znr3b U915 ( .A(FMREMNXT_7), .B(n2402), .C(n2401), .Y(EOF11263) );
    zoai2x4b U916 ( .A(n2457), .B(n2458), .C(n2459), .D(n2460), .E(n2461), .F(
        n2462), .G(n2463), .H(n2464), .Y(FRCHGCHKBIT) );
    zmux21lb U917 ( .A(n2483), .B(n2486), .S(INTTHRESHOLD[2]), .Y(n2457) );
    zor2b U918 ( .A(INTTHRESHOLD[5]), .B(n2509), .Y(n2459) );
    zivb U919 ( .A(INTTHRESHOLD[6]), .Y(n2511) );
    zor2b U920 ( .A(INTTHRESHOLD[7]), .B(INTTHRESHOLD[6]), .Y(n2462) );
    zxo2b U921 ( .A(n2496), .B(FRNUM[3]), .Y(n2464) );
    zivb U922 ( .A(FRNUMNXT_T_3), .Y(n2496) );
    zivb U923 ( .A(n2459), .Y(n2475) );
    zan2b U924 ( .A(RSTREMAIN_), .B(FMREMNXT_7), .Y(FMREMN1078_7) );
    zan2b U925 ( .A(CMDSTART), .B(TXSOF), .Y(CMDTXSOF1868) );
    zan3b U926 ( .A(sub_325_carry_1), .B(n2331), .C(RSTREMAIN_), .Y(
        FRAMECHG1090) );
    znr2b U927 ( .A(LTINT_PCLK), .B(n2444), .Y(LTINT_PCLK1831) );
    zivb U928 ( .A(LTINT), .Y(n2444) );
    zao21b U929 ( .A(SOFGEN), .B(FRCHGCHKBIT_2T), .C(GEN_PERR), .Y(LTINT) );
    zan2b U930 ( .A(RSTREMAIN_), .B(FMREMNXT_11), .Y(FMREMN1078_11) );
    zivb U931 ( .A(REDUCE), .Y(val313_4) );
    zan2b U932 ( .A(RSTREMAIN_), .B(FMREMNXT_5), .Y(FMREMN1078_5) );
    zan2b U933 ( .A(RSTREMAIN_), .B(FMREMNXT_2), .Y(FMREMN1078_2) );
    zoai21b U934 ( .A(n2440), .B(n2441), .C(n2442), .Y(ROLLCHKBIT) );
    zmux21lb U935 ( .A(n2517), .B(n2516), .S(FRLSTSIZE[1]), .Y(n2442) );
    zoai21b U936 ( .A(ASYNC_ACT), .B(n2446), .C(n2447), .Y(EHCIRESTART1600) );
    zmux21lb U937 ( .A(c1612_1), .B(b1610_1), .S(SLEEPTIME_SEL), .Y(n2447) );
    zan2b U938 ( .A(RSTREMAIN_), .B(FMREMNXT_3), .Y(FMREMN1078_3) );
    zan3b U939 ( .A(n1311), .B(RSTREMAIN_), .C(n1309), .Y(EOF21267) );
    znd3b U940 ( .A(n2425), .B(n2424), .C(n2423), .Y(n1311) );
    zan2b U941 ( .A(RSTREMAIN_), .B(FMREMNXT_10), .Y(FMREMN1078_10) );
    zan2b U942 ( .A(RSTREMAIN_), .B(FMREMNXT_4), .Y(FMREMN1078_4) );
    zivb U943 ( .A(n2450), .Y(RSTREMAIN_) );
    zor2b U944 ( .A(n2443), .B(WR_FRNUMT_T), .Y(FRNUM_PCLK_LATCH) );
    zivb U945 ( .A(FRNUM_PCLK_LATCH), .Y(n2519) );
    zivb U946 ( .A(FRLSTSIZE[1]), .Y(n2466) );
    zan2b U947 ( .A(FRNUM_PCLK[12]), .B(n2465), .Y(FRNUM_AD[12]) );
    zxo2b U948 ( .A(n2504), .B(FRLSTSIZE[1]), .Y(n2465) );
    zivb U949 ( .A(FRLSTSIZE[0]), .Y(n2504) );
    zivb U950 ( .A(n2465), .Y(n2441) );
    znr4b U951 ( .A(n2445), .B(CMDTXSOF_3T), .C(CMDTXSOF_T), .D(CMDTXSOF), .Y(
        EHCI_MAC_EOT) );
    zan2b U952 ( .A(ROLLOVER_S_T), .B(RUN), .Y(ROLLOVER_S) );
    zdffqrb FRNUM_W_reg_13 ( .CK(PCICLK), .D(FRNUM_W484_13), .R(TRST_), .Q(
        FRNUM_W_13) );
    zdffqrb FRNUM_W_reg_12 ( .CK(PCICLK), .D(FRNUM_W484_12), .R(TRST_), .Q(
        FRNUM_W_12) );
    zdffqrb FRNUM_W_reg_11 ( .CK(PCICLK), .D(FRNUM_W484_11), .R(TRST_), .Q(
        FRNUM_W_11) );
    zdffqrb FRNUM_W_reg_10 ( .CK(PCICLK), .D(FRNUM_W484_10), .R(TRST_), .Q(
        FRNUM_W_10) );
    zdffqrb FRNUM_W_reg_9 ( .CK(PCICLK), .D(FRNUM_W484_9), .R(TRST_), .Q(
        FRNUM_W_9) );
    zdffqrb FRNUM_W_reg_8 ( .CK(PCICLK), .D(FRNUM_W484_8), .R(TRST_), .Q(
        FRNUM_W_8) );
    zdffqrb FRNUM_W_reg_7 ( .CK(PCICLK), .D(FRNUM_W484_7), .R(TRST_), .Q(
        FRNUM_W_7) );
    zdffqrb FRNUM_W_reg_6 ( .CK(PCICLK), .D(FRNUM_W484_6), .R(TRST_), .Q(
        FRNUM_W_6) );
    zdffqrb FRNUM_W_reg_5 ( .CK(PCICLK), .D(FRNUM_W484_5), .R(TRST_), .Q(
        FRNUM_W_5) );
    zdffqrb FRNUM_W_reg_4 ( .CK(PCICLK), .D(FRNUM_W484_4), .R(TRST_), .Q(
        FRNUM_W_4) );
    zdffqrb FRNUM_W_reg_3 ( .CK(PCICLK), .D(FRNUM_W484_3), .R(TRST_), .Q(
        FRNUM_W_3) );
    zdffqrb FRNUM_W_reg_2 ( .CK(PCICLK), .D(FRNUM_W484_2), .R(TRST_), .Q(
        FRNUM_W_2) );
    zdffqrb FRNUM_W_reg_1 ( .CK(PCICLK), .D(FRNUM_W484_1), .R(TRST_), .Q(
        FRNUM_W_1) );
    zdffqrb FRNUM_W_reg_0 ( .CK(PCICLK), .D(FRNUM_W484_0), .R(TRST_), .Q(
        FRNUM_W_0) );
    zdffqrb FRNUM_PCLK_reg_13 ( .CK(PCICLK), .D(FRNUM_PCLK575_13), .R(TRST_), 
        .Q(FRNUM_PCLK[13]) );
    zdffqrb FRNUM_PCLK_reg_12 ( .CK(PCICLK), .D(FRNUM_PCLK575_12), .R(TRST_), 
        .Q(FRNUM_PCLK[12]) );
    zivb U953 ( .A(FRNUM_PCLK[12]), .Y(n2506) );
    zdffqrb FRNUM_PCLK_reg_11 ( .CK(PCICLK), .D(FRNUM_PCLK575_11), .R(TRST_), 
        .Q(FRNUM_PCLK[11]) );
    zivb U954 ( .A(FRNUM_PCLK[11]), .Y(n2507) );
    zdffqrb_ FRNUM_reg_13 ( .CK(CLK60M), .D(FRNUM730_13), .R(TRST_), .Q(FRNUM
        [13]) );
    zivb U955 ( .A(FRNUM[13]), .Y(n2440) );
    zdffqrb_ FRNUM_reg_12 ( .CK(CLK60M), .D(FRNUM730_12), .R(TRST_), .Q(FRNUM
        [12]) );
    zivb U956 ( .A(FRNUM[12]), .Y(n2499) );
    zdffqrb_ FRNUM_reg_11 ( .CK(CLK60M), .D(FRNUM730_11), .R(TRST_), .Q(FRNUM
        [11]) );
    zivb U957 ( .A(FRNUM[11]), .Y(n2500) );
    zdffqrb_ FRNUM_reg_10 ( .CK(CLK60M), .D(FRNUM730_10), .R(TRST_), .Q(FRNUM
        [10]) );
    zdffqrb_ FRNUM_reg_9 ( .CK(CLK60M), .D(FRNUM730_9), .R(TRST_), .Q(FRNUM[9]
        ) );
    zdffqrb_ FRNUM_reg_8 ( .CK(CLK60M), .D(FRNUM730_8), .R(TRST_), .Q(FRNUM[8]
        ) );
    zdffqrb_ FRNUM_reg_7 ( .CK(CLK60M), .D(FRNUM730_7), .R(TRST_), .Q(FRNUM[7]
        ) );
    zdffqrb_ FRNUM_reg_6 ( .CK(CLK60M), .D(FRNUM730_6), .R(TRST_), .Q(FRNUM[6]
        ) );
    zdffqrb_ FRNUM_reg_5 ( .CK(CLK60M), .D(FRNUM730_5), .R(TRST_), .Q(FRNUM[5]
        ) );
    zdffqrb_ FRNUM_reg_4 ( .CK(CLK60M), .D(FRNUM730_4), .R(TRST_), .Q(FRNUM[4]
        ) );
    zdffqrb_ FRNUM_reg_3 ( .CK(CLK60M), .D(FRNUM730_3), .R(TRST_), .Q(FRNUM[3]
        ) );
    zdffqrb_ FRNUM_reg_2 ( .CK(CLK60M), .D(FRNUM730_2), .R(TRST_), .Q(FRNUM[2]
        ) );
    zivb U958 ( .A(FRNUM[2]), .Y(n2469) );
    zdffqrb_ FRNUM_reg_1 ( .CK(CLK60M), .D(FRNUM730_1), .R(TRST_), .Q(FRNUM[1]
        ) );
    zivb U959 ( .A(FRNUM[1]), .Y(n2470) );
    zdffqrb_ SOFV_reg_10 ( .CK(CLK60M), .D(SOFV769_10), .R(TRST_), .Q(SOFV[10]
        ) );
    zdffqrb_ SOFV_reg_9 ( .CK(CLK60M), .D(SOFV769_9), .R(TRST_), .Q(SOFV[9])
         );
    zdffqrb_ SOFV_reg_8 ( .CK(CLK60M), .D(SOFV769_8), .R(TRST_), .Q(SOFV[8])
         );
    zdffqrb_ SOFV_reg_7 ( .CK(CLK60M), .D(SOFV769_7), .R(TRST_), .Q(SOFV[7])
         );
    zdffqrb_ SOFV_reg_6 ( .CK(CLK60M), .D(SOFV769_6), .R(TRST_), .Q(SOFV[6])
         );
    zdffqrb_ SOFV_reg_5 ( .CK(CLK60M), .D(SOFV769_5), .R(TRST_), .Q(SOFV[5])
         );
    zdffqrb_ SOFV_reg_4 ( .CK(CLK60M), .D(SOFV769_4), .R(TRST_), .Q(SOFV[4])
         );
    zdffqrb_ SOFV_reg_3 ( .CK(CLK60M), .D(SOFV769_3), .R(TRST_), .Q(SOFV[3])
         );
    zdffqrb_ SOFV_reg_2 ( .CK(CLK60M), .D(SOFV769_2), .R(TRST_), .Q(SOFV[2])
         );
    zdffqrb_ SOFV_reg_1 ( .CK(CLK60M), .D(SOFV769_1), .R(TRST_), .Q(SOFV[1])
         );
    zdffqrb_ SOFV_reg_0 ( .CK(CLK60M), .D(SOFV769_0), .R(TRST_), .Q(SOFV[0])
         );
    zdffqrb TMCNT_reg_12 ( .CK(CLK60M), .D(TMCNT1530_12), .R(TRST_), .Q(
        TMCNT_12) );
    zdffqrb TMCNT_reg_11 ( .CK(CLK60M), .D(TMCNT1530_11), .R(TRST_), .Q(
        TMCNT_11) );
    zdffqrb TMCNT_reg_10 ( .CK(CLK60M), .D(TMCNT1530_10), .R(TRST_), .Q(
        TMCNT_10) );
    zdffqrb TMCNT_reg_9 ( .CK(CLK60M), .D(TMCNT1530_9), .R(TRST_), .Q(TMCNT_9)
         );
    zdffqrb TMCNT_reg_8 ( .CK(CLK60M), .D(TMCNT1530_8), .R(TRST_), .Q(TMCNT_8)
         );
    zdffqrb TMCNT_reg_7 ( .CK(CLK60M), .D(TMCNT1530_7), .R(TRST_), .Q(TMCNT_7)
         );
    zdffqrb TMCNT_reg_6 ( .CK(CLK60M), .D(TMCNT1530_6), .R(TRST_), .Q(TMCNT_6)
         );
    zivb U960 ( .A(TMCNT_6), .Y(n2434) );
    zdffqrb TMCNT_reg_5 ( .CK(CLK60M), .D(TMCNT1530_5), .R(TRST_), .Q(TMCNT_5)
         );
    zdffqrb TMCNT_reg_4 ( .CK(CLK60M), .D(TMCNT1530_4), .R(TRST_), .Q(TMCNT_4)
         );
    zdffqrb TMCNT_reg_3 ( .CK(CLK60M), .D(TMCNT1530_3), .R(TRST_), .Q(TMCNT_3)
         );
    zdffqrb TMCNT_reg_2 ( .CK(CLK60M), .D(TMCNT1530_2), .R(TRST_), .Q(TMCNT_2)
         );
    zdffqrb TMCNT_reg_1 ( .CK(CLK60M), .D(TMCNT1530_1), .R(TRST_), .Q(TMCNT_1)
         );
    zdffqrb TMCNT_reg_0 ( .CK(CLK60M), .D(TMCNT1530_0), .R(TRST_), .Q(TMCNT_0)
         );
    zivb U961 ( .A(TMCNT_0), .Y(TMCNT1516_0) );
    zdffqrb HSERR_S_T_reg ( .CK(PCICLK), .D(HSERR_S), .R(TRST_), .Q(HSERR_S_T)
         );
    zdffqrb WR_FRNUMT_T_reg ( .CK(PCICLK), .D(WR_FRNUMT), .R(TRST_), .Q(
        WR_FRNUMT_T) );
    zdffqrb FMREMN_reg_12 ( .CK(CLK60M), .D(FMREMN1078_12), .R(TRST_), .Q(
        FMREMN_12) );
    zdffqrb FMREMN_reg_6 ( .CK(CLK60M), .D(FMREMN1078_6), .R(TRST_), .Q(
        FMREMN_6) );
    zdffqrb_ ROLLOVER_S_T_reg ( .CK(CLK60M), .D(n2525), .R(TRST_), .Q(
        ROLLOVER_S_T) );
    zdffqrb START_EVENT_T_reg ( .CK(PCICLK), .D(START_EVENT), .R(TRST_), .Q(
        START_EVENT_T) );
    zdffqsb FMREMN_reg_1 ( .CK(CLK60M), .D(FMREMN1078_1), .S(TRST_), .Q(
        FMREMN_1) );
    zivb U962 ( .A(FMREMN_1), .Y(n2503) );
    zdffqrb WR_FRNUMT_reg ( .CK(PCICLK), .D(WR_FRNUMT393), .R(TRST_), .Q(
        WR_FRNUMT) );
    zdffsb PRESOF_reg ( .CK(CLK60M), .D(PRESOF1203), .S(TRST_), .Q(PRESOF), 
        .QN(n2505) );
    zdffqrb_ HSERR_S_2T_reg ( .CK(PCICLK), .D(HSERR_S), .R(TRST_), .Q(
        HSERR_S_2T) );
    zdffqrb FMREMN_reg_8 ( .CK(CLK60M), .D(FMREMN1078_8), .R(TRST_), .Q(
        FMREMN_8) );
    zdffqrb ASYNCINT_reg ( .CK(LTINT_CK), .D(QHASYNCINT), .R(n2333), .Q(
        ASYNCINT) );
    zdffqrb START_EVENT_2T_reg ( .CK(PCICLK), .D(START_EVENT_T), .R(TRST_), 
        .Q(START_EVENT_2T) );
    zdffqrb TMCNT_EN_reg ( .CK(CLK60M), .D(TMCNT_EN1460), .R(TRST_), .Q(
        TMCNT_EN) );
    zivb U963 ( .A(TMCNT_EN), .Y(n2497) );
    zdffqrb FMREMN_reg_9 ( .CK(CLK60M), .D(FMREMN1078_9), .R(TRST_), .Q(
        FMREMN_9) );
    zdffqrb START_EVENT_SYNC_reg ( .CK(CLK60M), .D(START_EVENT_SYNC1423), .R(
        TRST_), .Q(START_EVENT_SYNC) );
    zdffqsb EOF1_reg ( .CK(CLK60M), .D(EOF11262), .S(TRST_), .Q(EOF1) );
    zdffqrb EHCI_MAC_EOT_PCLK_reg ( .CK(PCICLK), .D(MAC_EOT), .R(TRST_), .Q(
        EHCI_MAC_EOT_PCLK) );
    zdffqrb FRAMECHG_2T_reg ( .CK(PCICLK), .D(FRAMECHG_T), .R(TRST_), .Q(
        FRAMECHG_2T) );
    zdffqrb_ START_EVENT_3T_reg ( .CK(PCICLK), .D(START_EVENT_T), .R(TRST_), 
        .Q(START_EVENT_3T) );
    zdffqrb SOFGEN_reg ( .CK(CLK60M), .D(SOFGEN1084), .R(TRST_), .Q(SOFGEN) );
    zdffqrb_ FRCHGCHKBIT_T_reg ( .CK(CLK60M), .D(FRCHGCHKBIT), .R(TRST_), .Q(
        FRCHGCHKBIT_T) );
    zdffqrb FMREMN_reg_7 ( .CK(CLK60M), .D(FMREMN1078_7), .R(TRST_), .Q(
        FMREMN_7) );
    zdffqrb CMDTXSOF_reg ( .CK(PCICLK), .D(CMDTXSOF1868), .R(TRST_), .Q(
        CMDTXSOF) );
    zdffqrb FRAMECHG_reg ( .CK(CLK60M), .D(FRAMECHG1090), .R(TRST_), .Q(
        FRAMECHG) );
    zivb U964 ( .A(FRAMECHG), .Y(n2498) );
    zdffqrb FRAMECHG_T_reg ( .CK(PCICLK), .D(FRAMECHG), .R(TRST_), .Q(
        FRAMECHG_T) );
    zdffqrb LTINT_PCLK_reg ( .CK(PCICLK), .D(LTINT_PCLK1831), .R(TRST_), .Q(
        LTINT_PCLK) );
    zdffqrb CMDTXSOF_2T_reg ( .CK(PCICLK), .D(CMDTXSOF_T), .R(TRST_), .Q(
        CMDTXSOF_2T) );
    zdffqrb FMREMN_reg_11 ( .CK(CLK60M), .D(FMREMN1078_11), .R(TRST_), .Q(
        FMREMN_11) );
    zdffqrb FMREMN_reg_5 ( .CK(CLK60M), .D(FMREMN1078_5), .R(TRST_), .Q(
        FMREMN_5) );
    zdffqrb CMDTXSOF_3T_reg ( .CK(PCICLK), .D(CMDTXSOF_2T), .R(TRST_), .Q(
        CMDTXSOF_3T) );
    zdffqrb FMREMN_reg_2 ( .CK(CLK60M), .D(FMREMN1078_2), .R(TRST_), .Q(
        FMREMN_2) );
    zdffqrb_ ROLLCHKBIT_T_reg ( .CK(CLK60M), .D(ROLLCHKBIT), .R(TRST_), .Q(
        ROLLCHKBIT_T) );
    zdffqrb_ FRCHGCHKBIT_2T_reg ( .CK(CLK60M), .D(n2524), .R(TRST_), .Q(
        FRCHGCHKBIT_2T) );
    zdffrb EHCIRESTART_reg ( .CK(CLK60M), .D(EHCIRESTART1600), .R(TRST_), .Q(
        EHCIRESTART), .QN(n2446) );
    zdffqrb_ WR_FRNUMT_3T_reg ( .CK(PCICLK), .D(WR_FRNUMT), .R(TRST_), .Q(
        WR_FRNUMT_3T) );
    zdffqrb FMREMN_reg_3 ( .CK(CLK60M), .D(FMREMN1078_3), .R(TRST_), .Q(
        FMREMN_3) );
    zdffqrb CMDTXSOF_T_reg ( .CK(PCICLK), .D(CMDTXSOF), .R(TRST_), .Q(
        CMDTXSOF_T) );
    zdffqrb EOF2_reg ( .CK(CLK60M), .D(EOF21267), .R(TRST_), .Q(EOF2) );
    zdffqrb FMREMN_reg_10 ( .CK(CLK60M), .D(FMREMN1078_10), .R(TRST_), .Q(
        FMREMN_10) );
    zdffqrb WR_FRNUMT_2T_reg ( .CK(PCICLK), .D(WR_FRNUMT_T), .R(TRST_), .Q(
        WR_FRNUMT_2T) );
    zdffqrb FMREMN_reg_4 ( .CK(CLK60M), .D(FMREMN1078_4), .R(TRST_), .Q(
        FMREMN_4) );
    znr2d U965 ( .A(FROZSYNC), .B(n2514), .Y(n2326) );
    znr2b U966 ( .A(FROZSYNC), .B(n2497), .Y(n2327) );
    znr2d U967 ( .A(n2498), .B(n2451), .Y(n2328) );
    znr2d U968 ( .A(FRAMECHG), .B(n2451), .Y(n2329) );
    znr2b U969 ( .A(n2467), .B(n2451), .Y(n2330) );
    znr2b U970 ( .A(n2501), .B(n2503), .Y(n2331) );
    zivb U971 ( .A(FMREMNXT_7), .Y(n2423) );
    zivb U972 ( .A(FMREMNXT_6), .Y(n2406) );
    zivb U973 ( .A(FMREMNXT_9), .Y(n2409) );
    zivb U974 ( .A(FMREMNXT_10), .Y(n2410) );
    zivb U975 ( .A(FMREMNXT_6), .Y(n2424) );
    zivb U976 ( .A(FMREMNXT_4), .Y(n2419) );
    zivb U977 ( .A(FMREMNXT_2), .Y(n2412) );
    zivb U978 ( .A(FMREMNXT_3), .Y(n2396) );
    zivb U979 ( .A(FMREMNXT_5), .Y(n2399) );
    zivb U980 ( .A(FMREMNXT_11), .Y(n2403) );
    zxn2b U981 ( .A(MAXLEN[2]), .B(MAXLEN[0]), .Y(n2332) );
    zdffqrb_ FRNUM_reg_0 ( .CK(CLK60M), .D(FRNUM730_0), .R(TRST_), .Q(FRNUM[0]
        ) );
    zivb U982 ( .A(FRNUM[0]), .Y(n2468) );
    zor2b U983 ( .A(ATPG_ENI), .B(INTASYNC), .Y(n2333) );
    zdffqrb FMREMN_reg_0 ( .CK(CLK60M), .D(FMREMN1078_0), .R(TRST_), .Q(
        sub_325_carry_1) );
    zivb U984 ( .A(sub_325_carry_1), .Y(n2456) );
    zivb U985 ( .A(n2455), .Y(n2334) );
    zivb U986 ( .A(FROZSYNC), .Y(n2455) );
    zan2b U987 ( .A(FMREMN_10), .B(n2334), .Y(n2448) );
    zan2b U988 ( .A(FMREMN_8), .B(n2334), .Y(n2449) );
    zao22b U989 ( .A(n2334), .B(TMCNT_9), .C(n2327), .D(TMCNT1516_9), .Y(
        TMCNT1530_9) );
    zao22b U990 ( .A(TMCNT_12), .B(FROZSYNC), .C(TMCNT1516_12), .D(n2327), .Y(
        TMCNT1530_12) );
    zao22b U991 ( .A(TMCNT_3), .B(n2334), .C(TMCNT1516_3), .D(n2327), .Y(
        TMCNT1530_3) );
    zao22b U992 ( .A(TMCNT_11), .B(n2334), .C(TMCNT1516_11), .D(n2327), .Y(
        TMCNT1530_11) );
    zao22b U993 ( .A(TMCNT_5), .B(n2334), .C(TMCNT1516_5), .D(n2327), .Y(
        TMCNT1530_5) );
    zao22b U994 ( .A(TMCNT_1), .B(n2334), .C(TMCNT1516_1), .D(n2327), .Y(
        TMCNT1530_1) );
    zao22b U995 ( .A(TMCNT_6), .B(n2334), .C(TMCNT1516_6), .D(n2327), .Y(
        TMCNT1530_6) );
    zao22b U996 ( .A(TMCNT_0), .B(FROZSYNC), .C(TMCNT1516_0), .D(n2327), .Y(
        TMCNT1530_0) );
    zao22b U997 ( .A(TMCNT_4), .B(FROZSYNC), .C(TMCNT1516_4), .D(n2327), .Y(
        TMCNT1530_4) );
    zao22b U998 ( .A(TMCNT_8), .B(n2334), .C(TMCNT1516_8), .D(n2327), .Y(
        TMCNT1530_8) );
    zao22b U999 ( .A(TMCNT_2), .B(n2334), .C(TMCNT1516_2), .D(n2327), .Y(
        TMCNT1530_2) );
    zao22b U1000 ( .A(TMCNT_7), .B(n2334), .C(TMCNT1516_7), .D(n2327), .Y(
        TMCNT1530_7) );
    zao22b U1001 ( .A(TMCNT_10), .B(n2334), .C(TMCNT1516_10), .D(n2327), .Y(
        TMCNT1530_10) );
    zdffqsb FROZSYNC_reg ( .CK(CLK60M), .D(FROZEN), .S(TRST_), .Q(FROZSYNC) );
    zbfb U1002 ( .A(FRNUM_AD[0]), .Y(FRNUM_PCLK[0]) );
    zdffqrb FRNUM_PCLK_reg_0 ( .CK(PCICLK), .D(FRNUM_PCLK575_0), .R(TRST_), 
        .Q(FRNUM_AD[0]) );
    zbfb U1003 ( .A(FRNUM_AD[1]), .Y(FRNUM_PCLK[1]) );
    zdffqrb FRNUM_PCLK_reg_1 ( .CK(PCICLK), .D(FRNUM_PCLK575_1), .R(TRST_), 
        .Q(FRNUM_AD[1]) );
    zbfb U1004 ( .A(FRNUM_AD[2]), .Y(FRNUM_PCLK[2]) );
    zdffqrb FRNUM_PCLK_reg_2 ( .CK(PCICLK), .D(FRNUM_PCLK575_2), .R(TRST_), 
        .Q(FRNUM_AD[2]) );
    zbfb U1005 ( .A(FRNUM_AD[3]), .Y(FRNUM_PCLK[3]) );
    zdffqrb FRNUM_PCLK_reg_3 ( .CK(PCICLK), .D(FRNUM_PCLK575_3), .R(TRST_), 
        .Q(FRNUM_AD[3]) );
    zbfb U1006 ( .A(FRNUM_AD[4]), .Y(FRNUM_PCLK[4]) );
    zdffqrb FRNUM_PCLK_reg_4 ( .CK(PCICLK), .D(FRNUM_PCLK575_4), .R(TRST_), 
        .Q(FRNUM_AD[4]) );
    zbfb U1007 ( .A(FRNUM_AD[5]), .Y(FRNUM_PCLK[5]) );
    zdffqrb FRNUM_PCLK_reg_5 ( .CK(PCICLK), .D(FRNUM_PCLK575_5), .R(TRST_), 
        .Q(FRNUM_AD[5]) );
    zbfb U1008 ( .A(FRNUM_AD[6]), .Y(FRNUM_PCLK[6]) );
    zdffqrb FRNUM_PCLK_reg_6 ( .CK(PCICLK), .D(FRNUM_PCLK575_6), .R(TRST_), 
        .Q(FRNUM_AD[6]) );
    zbfb U1009 ( .A(FRNUM_AD[7]), .Y(FRNUM_PCLK[7]) );
    zdffqrb FRNUM_PCLK_reg_7 ( .CK(PCICLK), .D(FRNUM_PCLK575_7), .R(TRST_), 
        .Q(FRNUM_AD[7]) );
    zbfb U1010 ( .A(FRNUM_AD[8]), .Y(FRNUM_PCLK[8]) );
    zdffqrb FRNUM_PCLK_reg_8 ( .CK(PCICLK), .D(FRNUM_PCLK575_8), .R(TRST_), 
        .Q(FRNUM_AD[8]) );
    zbfb U1011 ( .A(FRNUM_AD[9]), .Y(FRNUM_PCLK[9]) );
    zdffqrb FRNUM_PCLK_reg_9 ( .CK(PCICLK), .D(FRNUM_PCLK575_9), .R(TRST_), 
        .Q(FRNUM_AD[9]) );
    zbfb U1012 ( .A(FRNUM_AD[10]), .Y(FRNUM_PCLK[10]) );
    zdffqrb FRNUM_PCLK_reg_10 ( .CK(PCICLK), .D(FRNUM_PCLK575_10), .R(TRST_), 
        .Q(FRNUM_AD[10]) );
    znr2b U1013 ( .A(n2377), .B(n2376), .Y(n2393) );
    zan2b U1014 ( .A(MAXLEN[10]), .B(add_378_carry_10), .Y(PRESOF_CAL_11) );
    zxo2b U1015 ( .A(MAXLEN[10]), .B(add_378_carry_10), .Y(PRESOF_CAL_10) );
    zan2b U1016 ( .A(MAXLEN[2]), .B(MAXLEN[0]), .Y(add_378_carry_1) );
    zan2b U1017 ( .A(add_378_2_carry_8), .B(MAXLEN[10]), .Y(n1131_23) );
    zxo2b U1018 ( .A(MAXLEN[10]), .B(add_378_2_carry_8), .Y(n1131_24) );
    zor2b U1019 ( .A(add_378_2_carry_7), .B(MAXLEN[9]), .Y(add_378_2_carry_8)
         );
    zxn2b U1020 ( .A(add_378_2_carry_7), .B(MAXLEN[9]), .Y(n1131_25) );
    zan2b U1021 ( .A(add_378_2_carry_6), .B(MAXLEN[8]), .Y(add_378_2_carry_7)
         );
    zxo2b U1022 ( .A(MAXLEN[8]), .B(add_378_2_carry_6), .Y(n1131_26) );
    zan2b U1023 ( .A(add_378_2_carry_5), .B(MAXLEN[7]), .Y(add_378_2_carry_6)
         );
    zxo2b U1024 ( .A(MAXLEN[7]), .B(add_378_2_carry_5), .Y(n1131_27) );
    zor2b U1025 ( .A(add_378_2_carry_4), .B(MAXLEN[6]), .Y(add_378_2_carry_5)
         );
    zxn2b U1026 ( .A(add_378_2_carry_4), .B(MAXLEN[6]), .Y(n1131_28) );
    zor2b U1027 ( .A(add_378_2_carry_3), .B(MAXLEN[5]), .Y(add_378_2_carry_4)
         );
    zxn2b U1028 ( .A(add_378_2_carry_3), .B(MAXLEN[5]), .Y(n1131_29) );
    zan2b U1029 ( .A(MAXLEN[3]), .B(MAXLEN[4]), .Y(add_378_2_carry_3) );
    zxo2b U1030 ( .A(MAXLEN[4]), .B(MAXLEN[3]), .Y(n1131_30) );
    zivb U1031 ( .A(MAXLEN[3]), .Y(n1131_31) );
    zan2b U1032 ( .A(FLADJ[4]), .B(add_60_carry_5), .Y(add_60_carry_6) );
    zxo2b U1033 ( .A(FLADJ[4]), .B(add_60_carry_5), .Y(FMINTV_5) );
    zan2b U1034 ( .A(FLADJ[3]), .B(add_60_carry_4), .Y(add_60_carry_5) );
    zxo2b U1035 ( .A(FLADJ[3]), .B(add_60_carry_4), .Y(FMINTV_4) );
    zan2b U1036 ( .A(FLADJ[0]), .B(REDUCE), .Y(add_60_carry_2) );
    zxo2b U1037 ( .A(FLADJ[0]), .B(REDUCE), .Y(FMINTV_1) );
    zfa1b add_60_U1_3 ( .A(val313_4), .B(FLADJ[2]), .CI(add_60_carry_3), .CO(
        add_60_carry_4), .S(FMINTV_3) );
    zfa1b add_60_U1_2 ( .A(val313_4), .B(FLADJ[1]), .CI(add_60_carry_2), .CO(
        add_60_carry_3), .S(FMINTV_2) );
    zfa1b add_60_U1_6 ( .A(REDUCE), .B(FLADJ[5]), .CI(add_60_carry_6), .CO(
        FMINTV_7), .S(FMINTV_6) );
    zfa1b add_378_U1_5 ( .A(MAXLEN[5]), .B(n1131_27), .CI(add_378_carry_5), 
        .CO(add_378_carry_6), .S(PRESOF_CAL_5) );
    zfa1b add_378_U1_4 ( .A(MAXLEN[4]), .B(n1131_28), .CI(add_378_carry_4), 
        .CO(add_378_carry_5), .S(PRESOF_CAL_4) );
    zfa1b add_378_U1_3 ( .A(MAXLEN[3]), .B(n1131_29), .CI(add_378_carry_3), 
        .CO(add_378_carry_4), .S(PRESOF_CAL_3) );
    zfa1b add_378_U1_9 ( .A(MAXLEN[9]), .B(n1131_23), .CI(add_378_carry_9), 
        .CO(add_378_carry_10), .S(PRESOF_CAL_9) );
    zfa1b add_378_U1_2 ( .A(MAXLEN[2]), .B(n1131_30), .CI(add_378_carry_2), 
        .CO(add_378_carry_3), .S(PRESOF_CAL_2) );
    zfa1b add_378_U1_7 ( .A(MAXLEN[7]), .B(n1131_25), .CI(add_378_carry_7), 
        .CO(add_378_carry_8), .S(PRESOF_CAL_7) );
    zfa1b add_378_U1_8 ( .A(MAXLEN[8]), .B(n1131_24), .CI(add_378_carry_8), 
        .CO(add_378_carry_9), .S(PRESOF_CAL_8) );
    zfa1b add_378_U1_6 ( .A(MAXLEN[6]), .B(n1131_26), .CI(add_378_carry_6), 
        .CO(add_378_carry_7), .S(PRESOF_CAL_6) );
    zfa1b add_378_U1_1 ( .A(MAXLEN[1]), .B(n1131_31), .CI(add_378_carry_1), 
        .CO(add_378_carry_2), .S(PRESOF_CAL_1) );
    zinr2b U1038 ( .A(n2399), .B(n2398), .Y(n2400) );
    zinr2b U1039 ( .A(n2423), .B(n2415), .Y(n1309) );
    zor3b U1040 ( .A(START_EVENT_2T), .B(START_EVENT_3T), .C(START_EVENT_T), 
        .Y(START_EVENT_SYNC1423) );
    zao222b U1041 ( .A(FMREMN_12), .B(FROZSYNC), .C(FMREMNXT957_12), .D(n2326), 
        .E(n2325), .F(val313_4), .Y(FMREMNXT_12) );
    zao222b U1042 ( .A(FMREMN_11), .B(FROZSYNC), .C(FMREMNXT957_11), .D(n2326), 
        .E(n2325), .F(val313_4), .Y(FMREMNXT_11) );
    zao211b U1043 ( .A(FMREMNXT957_10), .B(n2326), .C(n2325), .D(n2448), .Y(
        FMREMNXT_10) );
    zao222b U1044 ( .A(FMREMN_9), .B(FROZSYNC), .C(n2326), .D(FMREMNXT957_9), 
        .E(n2325), .F(REDUCE), .Y(FMREMNXT_9) );
    zao211b U1045 ( .A(FMREMNXT957_8), .B(n2326), .C(n2325), .D(n2449), .Y(
        FMREMNXT_8) );
    zao222b U1046 ( .A(FMREMN_7), .B(FROZSYNC), .C(FMREMNXT957_7), .D(n2326), 
        .E(FMINTV_7), .F(n2325), .Y(FMREMNXT_7) );
    zao222b U1047 ( .A(FMREMN_6), .B(FROZSYNC), .C(FMREMNXT957_6), .D(n2326), 
        .E(FMINTV_6), .F(n2325), .Y(FMREMNXT_6) );
    zao222b U1048 ( .A(FMREMN_5), .B(FROZSYNC), .C(FMREMNXT957_5), .D(n2326), 
        .E(FMINTV_5), .F(n2325), .Y(FMREMNXT_5) );
    zao222b U1049 ( .A(FMREMN_4), .B(FROZSYNC), .C(FMREMNXT957_4), .D(n2326), 
        .E(FMINTV_4), .F(n2325), .Y(FMREMNXT_4) );
    zao222b U1050 ( .A(FMREMN_3), .B(FROZSYNC), .C(FMREMNXT957_3), .D(n2326), 
        .E(FMINTV_3), .F(n2325), .Y(FMREMNXT_3) );
    zao222b U1051 ( .A(FMREMN_2), .B(FROZSYNC), .C(FMREMNXT957_2), .D(n2326), 
        .E(FMINTV_2), .F(n2325), .Y(FMREMNXT_2) );
    zao222b U1052 ( .A(FMREMN_1), .B(FROZSYNC), .C(FMREMNXT957_1), .D(n2326), 
        .E(FMINTV_1), .F(n2325), .Y(FMREMNXT_1) );
    zao222b U1053 ( .A(sub_325_carry_1), .B(FROZSYNC), .C(n2456), .D(n2326), 
        .E(REDUCE), .F(n2325), .Y(FMREMNXT_0) );
    zao222b U1054 ( .A(FRNUM_W_0), .B(n2451), .C(n2468), .D(n2328), .E(n2329), 
        .F(FRNUM[0]), .Y(FRNUM730_0) );
    zao222b U1055 ( .A(n2329), .B(FRNUM[1]), .C(FRNUM_W_1), .D(n2451), .E(
        FRNUMNXT_T_1), .F(n2328), .Y(FRNUM730_1) );
    zao222b U1056 ( .A(n2329), .B(FRNUM[2]), .C(FRNUM_W_2), .D(n2451), .E(
        FRNUMNXT_T_2), .F(n2328), .Y(FRNUM730_2) );
    zao222b U1057 ( .A(n2329), .B(FRNUM[3]), .C(FRNUM_W_3), .D(n2451), .E(
        FRNUMNXT_T_3), .F(n2328), .Y(FRNUM730_3) );
    zao222b U1058 ( .A(n2329), .B(FRNUM[4]), .C(FRNUM_W_4), .D(n2451), .E(
        FRNUMNXT_T_4), .F(n2328), .Y(FRNUM730_4) );
    zao222b U1059 ( .A(n2329), .B(FRNUM[5]), .C(FRNUM_W_5), .D(n2451), .E(
        FRNUMNXT_T_5), .F(n2328), .Y(FRNUM730_5) );
    zao222b U1060 ( .A(n2329), .B(FRNUM[6]), .C(FRNUM_W_6), .D(n2451), .E(
        FRNUMNXT_T_6), .F(n2328), .Y(FRNUM730_6) );
    zao222b U1061 ( .A(FRNUM_W_7), .B(n2451), .C(n2329), .D(FRNUM[7]), .E(
        FRNUMNXT_T_7), .F(n2328), .Y(FRNUM730_7) );
    zao222b U1062 ( .A(FRNUM_W_8), .B(n2451), .C(n2329), .D(FRNUM[8]), .E(
        FRNUMNXT_T_8), .F(n2328), .Y(FRNUM730_8) );
    zao222b U1063 ( .A(FRNUM_W_9), .B(n2451), .C(n2329), .D(FRNUM[9]), .E(
        n2328), .F(FRNUMNXT_T_9), .Y(FRNUM730_9) );
    zao222b U1064 ( .A(FRNUM_W_10), .B(n2451), .C(n2329), .D(FRNUM[10]), .E(
        FRNUMNXT_T_10), .F(n2328), .Y(FRNUM730_10) );
    zao222b U1065 ( .A(FRNUM_W_11), .B(n2451), .C(n2329), .D(FRNUM[11]), .E(
        FRNUMNXT_T_11), .F(n2328), .Y(FRNUM730_11) );
    zao222b U1066 ( .A(FRNUM_W_12), .B(n2451), .C(n2329), .D(FRNUM[12]), .E(
        FRNUMNXT_T_12), .F(n2328), .Y(FRNUM730_12) );
    zao222b U1067 ( .A(FRNUM_W_13), .B(n2451), .C(n2329), .D(FRNUM[13]), .E(
        FRNUMNXT_T_13), .F(n2328), .Y(FRNUM730_13) );
    zan4b U1068 ( .A(n2455), .B(n2456), .C(n2331), .D(RSTREMAIN_), .Y(
        SOFGEN1084) );
    zoa21d U1069 ( .A(FRLSTSIZE[0]), .B(n2466), .C(FRNUM_PCLK[11]), .Y(
        FRNUM_AD[11]) );
    zan4b U1070 ( .A(FRAMECHG), .B(n2468), .C(n2469), .D(n2470), .Y(n2467) );
    zinr2b U1071 ( .A(FRAMECHG_2T), .B(FRAMECHG_T), .Y(n2443) );
    zan4b U1072 ( .A(n2477), .B(n2478), .C(n2479), .D(n2480), .Y(n2463) );
    zoa21d U1073 ( .A(n2459), .B(n2481), .C(n2482), .Y(n2461) );
    zor3b U1074 ( .A(WR_FRNUMT_3T), .B(WR_FRNUMT), .C(WR_FRNUMT_T), .Y(n2451)
         );
    zor6b U1075 ( .A(FMREMN_6), .B(FMREMN_5), .C(FMREMN_4), .D(FMREMN_9), .E(
        FMREMN_11), .F(n2502), .Y(n2501) );
    zor4b U1076 ( .A(HSERR_S_T), .B(HSERR_S_2T), .C(HSERR_S), .D(n2471), .Y(
        n2450) );
    zor3b U1077 ( .A(FMREMN_1), .B(sub_325_carry_1), .C(n2501), .Y(n2515) );
    zor6b U1078 ( .A(FMREMN_12), .B(FMREMN_8), .C(FMREMN_3), .D(FMREMN_2), .E(
        FMREMN_7), .F(FMREMN_10), .Y(n2502) );
    zinr2b U1079 ( .A(EHCI_DBG_MAC_EOT), .B(SWDBG), .Y(n2472) );
    zor4b U1080 ( .A(INTTHRESHOLD[7]), .B(n2492), .C(n2510), .D(n2511), .Y(
        n2460) );
    zor3b U1081 ( .A(INTTHRESHOLD[5]), .B(n2510), .C(n2462), .Y(n2458) );
    zind2d U1082 ( .A(CMDTXSOF_2T), .B(EHCI_MAC_EOT_PCLK), .Y(n2445) );
    zor4b U1083 ( .A(n2510), .B(n2513), .C(n2494), .D(n2509), .Y(n2482) );
    zivb U1084 ( .A(FRCHGCHKBIT_T), .Y(n2523) );
    zivb U1085 ( .A(n2523), .Y(n2524) );
    zbfb U1086 ( .A(ROLLOVER_S_T633), .Y(n2525) );
endmodule


module AQHCTL ( QH_PARSE_GO, PARSEQHEND, QHPARSING, QHIDLE, DW0, DW1, DW2, DW3, 
    DW4, DW5, DW6, DW7, DW8, DW9, DW10, DW11, GEN_PERR, PCIEND, UP_DW3, UP_DW5, 
    UP_DW6, UP_DW7, UP_LDW3, UP_LDW5, UP_LDW6, UP_LDW7, CACHEPHASE, QHCIREQ, 
    QHDWNUM, QDWOFFSET, QHCIADR, QHCIADD, QHCIMWR, DWCNT, QHSM, TRAN_CMD, 
    QH_ACT, QBUI_GO, CACHE_ADDR, CACHE_INVALID, MAXLEN, CRCERR, ACTLEN, BABBLE, 
    PIDERR, TMOUT, RXNAK, RXNYET, RXSTALL, RXACK, RXDATA0, RXDATA1, RXPIDERR, 
    TOGMATCH, SPD, EHCI_MAC_EOT, FEMPTY, TDMAEND, QRXERR, QCMDSTART_REQ, 
    QCMDSTART, QEOT, QTDEXE, HEADSEEN, RECLAMATION, ASYNC_EMPTY, NAKCNTSM, 
    NAKCNTSMNXT, LTINT_PCLK, USBINT_EN, ERRINT_EN, USBINT, ERRINT, QHIOCINT_S, 
    QHERRINT_S, QHIOCINT, QHERRINT, PCICLK, EHCIFLOW_PCLK, TRST_ );
input  [31:0] DW0;
input  [31:0] DW1;
input  [31:0] DW6;
input  [31:0] DW7;
input  [31:0] DW9;
output [31:0] UP_DW6;
output [3:0] QDWOFFSET;
input  [1:0] NAKCNTSMNXT;
input  [26:0] CACHE_ADDR;
output [31:0] UP_DW7;
output [13:0] QHSM;
input  [1:0] NAKCNTSM;
input  [31:0] DW2;
input  [31:0] DW3;
input  [31:0] DW8;
input  [3:0] DWCNT;
input  [31:0] DW4;
output [31:0] UP_DW5;
output [31:0] QHCIADR;
output [31:0] QHCIADD;
input  [10:0] ACTLEN;
input  [31:0] DW5;
input  [31:0] DW10;
input  [31:0] DW11;
output [104:0] TRAN_CMD;
output [10:0] MAXLEN;
output [31:0] UP_DW3;
output [3:0] QHDWNUM;
input  QH_PARSE_GO, GEN_PERR, PCIEND, QH_ACT, CRCERR, BABBLE, PIDERR, TMOUT, 
    RXNAK, RXNYET, RXSTALL, RXACK, RXDATA0, RXDATA1, RXPIDERR, TOGMATCH, SPD, 
    EHCI_MAC_EOT, FEMPTY, TDMAEND, QCMDSTART, RECLAMATION, LTINT_PCLK, 
    USBINT_EN, ERRINT_EN, USBINT, ERRINT, PCICLK, EHCIFLOW_PCLK, TRST_;
output PARSEQHEND, QHPARSING, QHIDLE, UP_LDW3, UP_LDW5, UP_LDW6, UP_LDW7, 
    CACHEPHASE, QHCIREQ, QHCIMWR, QBUI_GO, CACHE_INVALID, QRXERR, 
    QCMDSTART_REQ, QEOT, QTDEXE, HEADSEEN, ASYNC_EMPTY, QHIOCINT_S, QHERRINT_S, 
    QHIOCINT, QHERRINT;
    wire VIR_TOTALBYTES_9, OVERWBOFFSET_P1671_9, OVERWBOFFSET1715_2, 
        VIR_TOTALBYTES_13, IMMEDRETRY1293, SPAREO6, MINUEND_8, TOTALBYTES640_7, 
        CERR1176_1, TOTALBYTES_12, TOTALBYTES_6, CURQTDPTR1422_20, 
        PARSEQHEND_PRE, NAKCNT1035_2, OVERWBOFFSET_P1671_0, VIR_TOTALBYTES_0, 
        QHERRINT2000, CURQTDPTR1422_15, QHSMNXT_12, NAKCNT996_3, 
        QHERRINT_T1963, TOTALBYTES640_14, CPAGE_0, CURQTDPTR1422_29, QHSMNXT_1, 
        TOTALBYTES_8, ASYNC_EMPTY1852, QHIOCINT_T1889, MINUEND_6, 
        TOTALBYTES640_13, SPAREO0_, TOTALBYTES640_9, CPAGE1098_0, SPAREO8, 
        CURQTDPTR1422_12, VIR_TOTALBYTES_7, OVERWBOFFSET_P1671_7, MINUEND_10, 
        TOTALBYTES_1, OVERWBOFFSET_P1671_11, CURQTDPTR1422_27, XACTERR1233, 
        CPAGE1102_2, TOTALBYTES640_0, VIR_TOTALBYTES_14, SPAREO1, 
        OVERWBOFFSET1715_5, CURQTDPTR1422_13, OVERWBOFFSET_P1671_6, 
        VIR_TOTALBYTES_6, CPAGE1098_1, SPAREO9, QCMDSTART_EOT, 
        PHASENXT_resultwb, MINUEND_7, TOTALBYTES640_12, TOTALBYTES640_8, 
        PHASENXT_idle, IMMEDRETRY, TOTALBYTES_9, QHSMNXT_7, CURQTDPTR1422_5, 
        OVERWBOFFSET1715_4, SPAREO0, TOTALBYTES640_1, TOTALBYTES_0, 
        OVERWBOFFSET_P1671_10, CURQTDPTR1422_26, TOTALBYTES_14, CERR1176_0, 
        QEOT1815, TOTALBYTES_7, TOTALBYTES_13, CURQTDPTR1422_21, n3187, 
        MINUEND_9, TOTALBYTES640_6, PING_ERR783, VIR_TOTALBYTES_12, SPAREO7, 
        SPLITXSTATE1256, OVERWBOFFSET_P1671_8, VIR_TOTALBYTES_8, 
        OVERWBOFFSET1715_3, CPAGE_1, CURQTDPTR1422_28, QHSMNXT_13, NAKCNT996_2, 
        NAKCNT1035_3, VIR_TOTALBYTES_1, OVERWBOFFSET_P1671_1, CURQTDPTR1422_14, 
        OVERWBOFFSET1715_1, ACTIVE, ACTIVE_NXT, QTDHALT, SPAREO5, 
        VIR_TOTALBYTES_10, TOTALBYTES640_4, TOTALBYTES_11, CURQTDPTR1422_23, 
        TOTALBYTES_5, LENGTMAX, OVERWBOFFSET1715_8, CURQTDPTR1422_9, 
        CURQTDPTR1422_16, NAKCNT1035_1, OVERWBOFFSET_P1671_3, CURQTDPTR1422_31, 
        VIR_TOTALBYTES_3, NAKCNT996_0, QHSMNXT_2, QHSMNXT_5, TOTALBYTES640_10, 
        MINUEND_5, QHIOCINT_T, DT881, ACCEPT_DATA, VIR_TOTALBYTES_4, 
        OVERWBOFFSET_P1671_4, OVERWBOFFSET1715_10, CURQTDPTR1422_11, 
        CURQTDPTR1422_24, OVERWBOFFSET_P1671_12, TOTALBYTES_2, CACHE_MODIFY497, 
        CERR_1, TOTALBYTES640_3, CPAGE1102_1, PING_PRESERVE, SPAREO2, 
        OVERWBOFFSET1715_6, CURQTDPTR1422_7, CURQTDPTR1422_18, 
        OVERWBOFFSET_P1671_5, VIR_TOTALBYTES_5, OVERWBOFFSET1715_11, 
        CURQTDPTR1422_10, CPAGE1098_2, TOTALBYTES640_11, MINUEND_4, QHSMNXT_4, 
        OVERWBOFFSET1715_7, CURQTDPTR1422_6, CURQTDPTR1422_19, QRXERR_CUR1331, 
        SPAREO3, QHIOCINT1926, SPAREO1_, CERR1180_1, CERR_0, TOTALBYTES640_2, 
        CACHE_INVALID1602, CURQTDPTR1422_25, QCMDSTART_EOT1778, CACHE_MODIFY, 
        TOTALBYTES_3, TOTALBYTES_10, CURQTDPTR1422_22, TOTALBYTES_4, 
        TOTALBYTES640_5, SPAREO4, VIR_TOTALBYTES_11, OVERWBOFFSET1715_0, 
        QHERRINT_T, CPAGE_2, PHASENXT_exechk, MINUEND_3, NAKCNT996_1, 
        QHSMNXT_10, OVERWBOFFSET1715_9, CURQTDPTR1422_8, CURQTDPTR1422_17, 
        NAKCNT1035_0, CURQTDPTR1422_30, VIR_TOTALBYTES_2, OVERWBOFFSET_P1671_2, 
        n2069, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
        n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2314, 
        n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, 
        n2325, n2326, n2327, n2328, n2358, n2428, n2429, n2430, n2431, n2432, 
        n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
        n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
        n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
        n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
        n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
        n2483, n2484, n2485, n2486, n2487, n2488, n2489, add_503_carry_2, 
        sub_383_carry_1, sub_383_B_not_10, sub_383_B_not_8, sub_383_carry_8, 
        sub_383_B_not_6, sub_383_carry_14, sub_383_carry_13, sub_383_carry_12, 
        sub_383_carry_7, sub_383_carry_6, sub_383_B_not_7, sub_383_B_not_9, 
        sub_383_carry_9, sub_383_carry_2, sub_383_B_not_5, sub_383_carry_11, 
        sub_383_carry_10, sub_383_carry_5, sub_383_carry_4, sub_383_B_not_4, 
        sub_383_carry_3, sub_383_B_not_3, n2490, r285_carry_8, r285_carry_1, 
        r285_carry_7, r285_carry_6, r285_carry_9, r285_carry_2, r285_carry_11, 
        r285_carry_10, r285_carry_5, r285_carry_4, r285_carry_3, n2491, n2492, 
        n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
        n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
        n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
        n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, 
        n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, 
        n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, 
        n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, 
        n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, 
        n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, 
        n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, 
        n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, 
        n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, 
        n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, 
        n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
        n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, 
        n2643, n2644, n2645, n2646, n2647, n2648, n2650, n2651, n2652, n2653, 
        n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, 
        n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, 
        n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, 
        n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, 
        n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, 
        n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, 
        n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, 
        n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, 
        n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, 
        n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, 
        n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, 
        n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, 
        n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, 
        n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
        n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, 
        n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, 
        n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, 
        n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, 
        n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, 
        n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, 
        n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, 
        n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, 
        n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, 
        n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, 
        n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, 
        n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, 
        n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, 
        n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, 
        n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, 
        n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, 
        n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
        n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
        n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
        n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
        n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, 
        n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
        n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
        n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
        n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
        n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
        n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
        n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
        n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
        n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
        n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
        n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
        n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
        n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
        n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
        n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
        n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
        n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, 
        n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
        n3184, n3185, n3186, _cell_705_U89_Z_10, _cell_705_U89_Z_9, 
        _cell_705_U89_Z_8, _cell_705_U89_Z_7, _cell_705_U89_Z_6, 
        _cell_705_U89_Z_5, _cell_705_U89_Z_4, _cell_705_U89_Z_3, 
        _cell_705_U89_Z_2, _cell_705_U89_Z_1, _cell_705_U89_Z_0;
    assign UP_DW3[4] = 1'b0;
    assign UP_DW3[3] = 1'b0;
    assign UP_DW3[2] = 1'b0;
    assign UP_DW3[1] = 1'b0;
    assign UP_DW3[0] = 1'b0;
    assign QDWOFFSET[3] = 1'b0;
    assign QDWOFFSET[2] = 1'b1;
    assign QDWOFFSET[1] = 1'b0;
    assign QDWOFFSET[0] = 1'b0;
    assign QHCIADR[4] = 1'b0;
    assign QHCIADR[1] = 1'b0;
    assign QHCIADR[0] = 1'b0;
    assign TRAN_CMD[51] = 1'b0;
    assign TRAN_CMD[12] = 1'b0;
    assign TRAN_CMD[10] = 1'b0;
    assign TRAN_CMD[2] = 1'b0;
    assign TRAN_CMD[1] = 1'b0;
    assign TRAN_CMD[0] = 1'b0;
    zoai21b SPARE845 ( .A(SPAREO1), .B(n2321), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE842 ( .A(SPAREO0), .B(n2319), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zaoi211b SPARE843 ( .A(SPAREO4), .B(PARSEQHEND_PRE), .C(SPAREO6), .D(1'b0), 
        .Y(SPAREO8) );
    zoai21b SPARE844 ( .A(SPAREO0), .B(SPAREO8), .C(ACCEPT_DATA), .Y(SPAREO9)
         );
    znr3b SPARE846 ( .A(SPAREO2), .B(LENGTMAX), .C(SPAREO0_), .Y(SPAREO4) );
    zdffrb SPARE841 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE848 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE840 ( .CK(PCICLK), .D(PING_PRESERVE), .R(1'b1), .Q(SPAREO0), 
        .QN(SPAREO0_) );
    znd3b SPARE849 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb SPARE847 ( .A(SPAREO4), .Y(SPAREO5) );
    znd2b U761 ( .A(TOTALBYTES_1), .B(n2480), .Y(n2447) );
    znd2b U762 ( .A(TOTALBYTES_2), .B(n2454), .Y(n2448) );
    zivb U763 ( .A(DW1[18]), .Y(n2454) );
    znd2b U764 ( .A(TOTALBYTES_0), .B(n2449), .Y(n2478) );
    zivb U765 ( .A(DW1[16]), .Y(n2449) );
    znr2b U766 ( .A(TOTALBYTES_1), .B(n2480), .Y(n2481) );
    zivb U767 ( .A(DW1[17]), .Y(n2480) );
    znd2b U768 ( .A(TOTALBYTES_3), .B(n2453), .Y(n2443) );
    zivb U769 ( .A(DW1[19]), .Y(n2453) );
    znd2b U770 ( .A(TOTALBYTES_4), .B(n2455), .Y(n2444) );
    zivb U771 ( .A(DW1[20]), .Y(n2455) );
    znd2b U772 ( .A(n2446), .B(n2445), .Y(n2474) );
    znd2b U773 ( .A(DW1[19]), .B(n3004), .Y(n2446) );
    znd2b U774 ( .A(DW1[18]), .B(n3006), .Y(n2445) );
    znr2b U775 ( .A(n2479), .B(n2476), .Y(n2477) );
    znr2b U776 ( .A(n2481), .B(n2478), .Y(n2479) );
    znd2b U777 ( .A(n2448), .B(n2447), .Y(n2476) );
    znd2b U778 ( .A(TOTALBYTES_5), .B(n2452), .Y(n2439) );
    zivb U779 ( .A(DW1[21]), .Y(n2452) );
    znd2b U780 ( .A(TOTALBYTES_6), .B(n2456), .Y(n2440) );
    zivb U781 ( .A(DW1[22]), .Y(n2456) );
    znd2b U782 ( .A(n2442), .B(n2441), .Y(n2470) );
    znd2b U783 ( .A(DW1[21]), .B(n3000), .Y(n2442) );
    znd2b U784 ( .A(DW1[20]), .B(n3002), .Y(n2441) );
    znr2b U785 ( .A(n2475), .B(n2472), .Y(n2473) );
    znr2b U786 ( .A(n2477), .B(n2474), .Y(n2475) );
    znd2b U787 ( .A(n2444), .B(n2443), .Y(n2472) );
    znd2b U788 ( .A(TOTALBYTES_7), .B(n2451), .Y(n2435) );
    zivb U789 ( .A(DW1[23]), .Y(n2451) );
    znd2b U790 ( .A(TOTALBYTES_8), .B(n2457), .Y(n2436) );
    zivb U791 ( .A(DW1[24]), .Y(n2457) );
    znd2b U792 ( .A(n2438), .B(n2437), .Y(n2466) );
    znd2b U793 ( .A(DW1[23]), .B(n2996), .Y(n2438) );
    znd2b U794 ( .A(DW1[22]), .B(n2998), .Y(n2437) );
    znr2b U795 ( .A(n2471), .B(n2468), .Y(n2469) );
    znr2b U796 ( .A(n2473), .B(n2470), .Y(n2471) );
    znd2b U797 ( .A(n2440), .B(n2439), .Y(n2468) );
    znd2b U798 ( .A(TOTALBYTES_10), .B(n2458), .Y(n2431) );
    znd2b U799 ( .A(TOTALBYTES_9), .B(n2450), .Y(n2432) );
    zivb U800 ( .A(DW1[25]), .Y(n2450) );
    znd2b U801 ( .A(n2434), .B(n2433), .Y(n2462) );
    znd2b U802 ( .A(DW1[25]), .B(n2992), .Y(n2434) );
    znd2b U803 ( .A(DW1[24]), .B(n2994), .Y(n2433) );
    znr2b U804 ( .A(n2467), .B(n2464), .Y(n2465) );
    znr2b U805 ( .A(n2469), .B(n2466), .Y(n2467) );
    znd2b U806 ( .A(n2436), .B(n2435), .Y(n2464) );
    zoai211b U807 ( .A(RXDATA1), .B(RXDATA0), .C(TOGMATCH), .D(TRAN_CMD[9]), 
        .Y(n2904) );
    zoai21b U808 ( .A(n3135), .B(VIR_TOTALBYTES_14), .C(n3139), .Y(n2962) );
    znd8b U809 ( .A(n3035), .B(n3136), .C(n3041), .D(n3040), .E(n3043), .F(
        n3028), .G(n3134), .H(n3038), .Y(n3135) );
    znd8b U810 ( .A(n2993), .B(n2999), .C(n2997), .D(n3003), .E(n3001), .F(
        n3005), .G(n3007), .H(n3009), .Y(n2919) );
    zan3b U811 ( .A(RXNAK), .B(n2896), .C(TRAN_CMD[7]), .Y(n2895) );
    znr2b U812 ( .A(TOTALBYTES_10), .B(n2458), .Y(n2459) );
    zivb U813 ( .A(DW1[26]), .Y(n2458) );
    znr2b U814 ( .A(n2463), .B(n2460), .Y(n2461) );
    znr2b U815 ( .A(n2465), .B(n2462), .Y(n2463) );
    znd2b U816 ( .A(n2432), .B(n2431), .Y(n2460) );
    znd2b U817 ( .A(n2429), .B(n2428), .Y(n2430) );
    zor2b U818 ( .A(RXNAK), .B(RXNYET), .Y(n2979) );
    zor2b U819 ( .A(QHSM[9]), .B(QHCIMWR), .Y(n2921) );
    zor2b U820 ( .A(n2508), .B(n2963), .Y(n2964) );
    zoai2x4b U821 ( .A(n2974), .B(n3055), .C(n3047), .D(n3048), .E(n3113), .F(
        n3114), .G(n3115), .H(n3116), .Y(n3112) );
    zivb U822 ( .A(n2965), .Y(n3115) );
    zivb U823 ( .A(n2964), .Y(n3116) );
    zan2b U824 ( .A(n2292), .B(n2502), .Y(n2924) );
    zmux21lb U825 ( .A(CERR_1), .B(CERR1180_1), .S(n3153), .Y(n2952) );
    zxo2b U826 ( .A(n2490), .B(CERR_0), .Y(CERR1180_1) );
    zao21b U827 ( .A(n2490), .B(n3045), .C(n2899), .Y(n3044) );
    zmux21lb U828 ( .A(CERR_0), .B(n3045), .S(n3153), .Y(n2955) );
    zivb U829 ( .A(n3046), .Y(n3153) );
    zor2b U830 ( .A(n2900), .B(n3044), .Y(n3046) );
    zmux21hb U831 ( .A(MAXLEN[0]), .B(ACTLEN[0]), .S(UP_DW6[8]), .Y(
        _cell_705_U89_Z_0) );
    zmux21hb U832 ( .A(MAXLEN[1]), .B(ACTLEN[1]), .S(TRAN_CMD[9]), .Y(
        _cell_705_U89_Z_1) );
    zmux21hb U833 ( .A(MAXLEN[2]), .B(ACTLEN[2]), .S(UP_DW6[8]), .Y(
        _cell_705_U89_Z_2) );
    zmux21hb U834 ( .A(MAXLEN[3]), .B(ACTLEN[3]), .S(TRAN_CMD[9]), .Y(
        _cell_705_U89_Z_3) );
    zmux21hb U835 ( .A(MAXLEN[4]), .B(ACTLEN[4]), .S(UP_DW6[8]), .Y(
        _cell_705_U89_Z_4) );
    zmux21hb U836 ( .A(MAXLEN[5]), .B(ACTLEN[5]), .S(TRAN_CMD[9]), .Y(
        _cell_705_U89_Z_5) );
    zmux21hb U837 ( .A(MAXLEN[6]), .B(ACTLEN[6]), .S(UP_DW6[8]), .Y(
        _cell_705_U89_Z_6) );
    zmux21hb U838 ( .A(MAXLEN[7]), .B(ACTLEN[7]), .S(TRAN_CMD[9]), .Y(
        _cell_705_U89_Z_7) );
    zmux21hb U839 ( .A(MAXLEN[8]), .B(ACTLEN[8]), .S(UP_DW6[8]), .Y(
        _cell_705_U89_Z_8) );
    zmux21hb U840 ( .A(MAXLEN[9]), .B(ACTLEN[9]), .S(UP_DW6[8]), .Y(
        _cell_705_U89_Z_9) );
    zmux21hb U841 ( .A(MAXLEN[10]), .B(ACTLEN[10]), .S(TRAN_CMD[9]), .Y(
        _cell_705_U89_Z_10) );
    zan3b U842 ( .A(n2904), .B(n2905), .C(n2906), .Y(n2903) );
    zivb U843 ( .A(n2319), .Y(n3139) );
    zao21b U844 ( .A(TRAN_CMD[14]), .B(TRAN_CMD[9]), .C(n2515), .Y(n2069) );
    znd2b U845 ( .A(n2484), .B(n2483), .Y(n2485) );
    znd2b U846 ( .A(UP_DW5[2]), .B(UP_DW5[1]), .Y(n2488) );
    znd2b U847 ( .A(n2487), .B(NAKCNT996_0), .Y(n2489) );
    zmux21lb U848 ( .A(RXNAK), .B(RXNYET), .S(n2524), .Y(n3085) );
    zan2b U849 ( .A(RXACK), .B(n2521), .Y(n2948) );
    znd4b U850 ( .A(n3093), .B(n3094), .C(n3030), .D(OVERWBOFFSET_P1671_12), 
        .Y(n3092) );
    zivb U851 ( .A(n3080), .Y(n3093) );
    zor2b U852 ( .A(TRAN_CMD[5]), .B(n3024), .Y(n3080) );
    zor2b U853 ( .A(QHSM[1]), .B(n3089), .Y(n3088) );
    zivb U854 ( .A(RXACK), .Y(n2905) );
    zan3b U855 ( .A(n2521), .B(TRAN_CMD[6]), .C(n2908), .Y(n2907) );
    zao32b U856 ( .A(n3138), .B(n2980), .C(n2900), .D(RXNAK), .E(TRAN_CMD[7]), 
        .Y(n2908) );
    zivb U857 ( .A(RXSTALL), .Y(n3138) );
    zivb U858 ( .A(RXNYET), .Y(n2980) );
    zivb U859 ( .A(RXNAK), .Y(n2961) );
    zan2b U860 ( .A(PING_PRESERVE), .B(n2521), .Y(n2520) );
    zoai21b U861 ( .A(n2660), .B(n3098), .C(n3104), .Y(n3100) );
    zmux21lb U862 ( .A(n3099), .B(RXACK), .S(UP_DW6[0]), .Y(n3098) );
    zivb U863 ( .A(n2979), .Y(n3099) );
    zoa22b U864 ( .A(n2937), .B(n2938), .C(n2939), .D(n2662), .Y(n2936) );
    zivb U865 ( .A(RXPIDERR), .Y(n2937) );
    zor2b U866 ( .A(n2899), .B(n2662), .Y(n2938) );
    zao22b U867 ( .A(TRAN_CMD[5]), .B(n2534), .C(DW6[0]), .D(n2943), .Y(n2941)
         );
    zor2b U868 ( .A(n2918), .B(DW5[0]), .Y(n3087) );
    znr8b U869 ( .A(n2919), .B(DW6[29]), .C(DW6[27]), .D(DW6[30]), .E(DW6[23]), 
        .F(DW6[26]), .G(DW6[25]), .H(DW6[28]), .Y(n2918) );
    zoa211b U870 ( .A(QHSM[6]), .B(QHSM[8]), .C(QH_ACT), .D(EHCI_MAC_EOT), .Y(
        n3023) );
    zan2b U871 ( .A(RXPIDERR), .B(TRAN_CMD[5]), .Y(n2897) );
    zoa22b U872 ( .A(n2302), .B(n2891), .C(FEMPTY), .D(n2892), .Y(n2890) );
    zivb U873 ( .A(DW6[15]), .Y(n3062) );
    zivb U874 ( .A(n2892), .Y(n3146) );
    zivb U875 ( .A(n2971), .Y(n3145) );
    zor2b U876 ( .A(QRXERR), .B(BABBLE), .Y(n3150) );
    zao21b U877 ( .A(QHSMNXT_10), .B(n2977), .C(n2893), .Y(n2521) );
    zao32b U878 ( .A(n2950), .B(n2534), .C(n2940), .D(n3104), .E(n3106), .Y(
        n3105) );
    zor2b U879 ( .A(TRAN_CMD[5]), .B(n3026), .Y(n3106) );
    zan3b U880 ( .A(n3104), .B(n2511), .C(n3030), .Y(n3103) );
    zor2b U881 ( .A(n2899), .B(n3024), .Y(n3026) );
    zor2b U882 ( .A(n2942), .B(n2501), .Y(n2949) );
    zoa22b U883 ( .A(n2512), .B(n2916), .C(n2497), .D(n2917), .Y(n2915) );
    zivb U884 ( .A(n2916), .Y(n3144) );
    zor2b U885 ( .A(n3084), .B(n3050), .Y(n3154) );
    zivb U886 ( .A(n3132), .Y(n3084) );
    zivb U887 ( .A(n3054), .Y(n3143) );
    zoa22b U888 ( .A(n2512), .B(n2913), .C(n2914), .D(n2497), .Y(n2912) );
    zor2b U889 ( .A(QHSM[6]), .B(QHSM[5]), .Y(n2963) );
    zor2b U890 ( .A(n2965), .B(n2972), .Y(n2973) );
    zivb U891 ( .A(n2963), .Y(n3113) );
    znr6b U892 ( .A(n2934), .B(MAXLEN[1]), .C(MAXLEN[0]), .D(MAXLEN[2]), .E(
        MAXLEN[4]), .F(MAXLEN[3]), .Y(n2933) );
    znr3b U893 ( .A(n2430), .B(TOTALBYTES_14), .C(TOTALBYTES_13), .Y(n2482) );
    zor2b U894 ( .A(TRAN_CMD[14]), .B(n2515), .Y(n2896) );
    zor2b U895 ( .A(n3071), .B(n3072), .Y(n3075) );
    zivb U896 ( .A(DWCNT[3]), .Y(n3071) );
    zivb U897 ( .A(n3066), .Y(n3147) );
    zor2b U898 ( .A(DWCNT[3]), .B(n3065), .Y(n3066) );
    zivb U899 ( .A(DWCNT[0]), .Y(n3065) );
    zor2b U900 ( .A(QHDWNUM[0]), .B(n3067), .Y(n3068) );
    zivb U901 ( .A(n3073), .Y(n3141) );
    zor2b U902 ( .A(DWCNT[3]), .B(n3072), .Y(n3073) );
    zivb U903 ( .A(n3069), .Y(n3149) );
    zor2b U904 ( .A(DWCNT[0]), .B(DWCNT[3]), .Y(n3069) );
    zivb U905 ( .A(n3067), .Y(n3142) );
    zoai2x4b U906 ( .A(n2650), .B(n3049), .C(n3121), .D(n2942), .E(n2888), .F(
        n2889), .G(CACHE_MODIFY), .H(n3122), .Y(n2494) );
    zivb U907 ( .A(n2966), .Y(n3121) );
    zor2b U908 ( .A(n2964), .B(n2965), .Y(n2966) );
    zivb U909 ( .A(n2927), .Y(n2888) );
    zivb U910 ( .A(n2926), .Y(n2889) );
    zor2b U911 ( .A(QHSM[1]), .B(n2966), .Y(n2926) );
    zivb U912 ( .A(n2972), .Y(n3118) );
    zan2b U913 ( .A(n2923), .B(n2502), .Y(n2922) );
    zmux21lb U914 ( .A(n2296), .B(n2958), .S(PCIEND), .Y(n3097) );
    zan2b U915 ( .A(n2295), .B(n2959), .Y(n2958) );
    zao32b U916 ( .A(n3083), .B(n2293), .C(n3132), .D(n2302), .E(n3148), .Y(
        n3155) );
    zivb U917 ( .A(n3050), .Y(n3083) );
    zivb U918 ( .A(n2891), .Y(n3148) );
    zivb U919 ( .A(n3155), .Y(n3122) );
    zivb U920 ( .A(VIR_TOTALBYTES_12), .Y(n3039) );
    zivb U921 ( .A(VIR_TOTALBYTES_11), .Y(n3040) );
    zmux21lb U922 ( .A(n3017), .B(n2951), .S(n2320), .Y(CERR1176_1) );
    zan2b U923 ( .A(n2952), .B(n2953), .Y(n2951) );
    zmux21lb U924 ( .A(n3018), .B(n2954), .S(n2320), .Y(CERR1176_0) );
    zan2b U925 ( .A(n2955), .B(n2953), .Y(n2954) );
    zivb U926 ( .A(VIR_TOTALBYTES_2), .Y(n3037) );
    zivb U927 ( .A(MINUEND_4), .Y(sub_383_B_not_4) );
    zivb U928 ( .A(VIR_TOTALBYTES_4), .Y(n3035) );
    zivb U929 ( .A(MINUEND_3), .Y(sub_383_B_not_3) );
    zivb U930 ( .A(VIR_TOTALBYTES_3), .Y(n3036) );
    zivb U931 ( .A(MINUEND_6), .Y(sub_383_B_not_6) );
    zivb U932 ( .A(VIR_TOTALBYTES_6), .Y(n3033) );
    zivb U933 ( .A(MINUEND_5), .Y(sub_383_B_not_5) );
    zivb U934 ( .A(VIR_TOTALBYTES_5), .Y(n3034) );
    zivb U935 ( .A(MINUEND_8), .Y(sub_383_B_not_8) );
    zivb U936 ( .A(VIR_TOTALBYTES_8), .Y(n3031) );
    zivb U937 ( .A(MINUEND_7), .Y(sub_383_B_not_7) );
    zivb U938 ( .A(VIR_TOTALBYTES_7), .Y(n3032) );
    zivb U939 ( .A(MINUEND_9), .Y(sub_383_B_not_9) );
    zivb U940 ( .A(VIR_TOTALBYTES_9), .Y(n3028) );
    zxo2b U941 ( .A(add_503_carry_2), .B(n2328), .Y(CPAGE1102_2) );
    zivb U942 ( .A(n2938), .Y(n3140) );
    zivb U943 ( .A(n3024), .Y(ACCEPT_DATA) );
    zor2b U944 ( .A(n2938), .B(n3080), .Y(n3081) );
    zivb U945 ( .A(VIR_TOTALBYTES_13), .Y(n3038) );
    zivb U946 ( .A(MINUEND_10), .Y(sub_383_B_not_10) );
    zivb U947 ( .A(VIR_TOTALBYTES_10), .Y(n3041) );
    zivb U948 ( .A(VIR_TOTALBYTES_1), .Y(n3042) );
    zivd U949 ( .A(n3029), .Y(n2663) );
    zivd U950 ( .A(n3027), .Y(n2664) );
    zor2b U951 ( .A(n2319), .B(n3026), .Y(n3027) );
    zivb U952 ( .A(VIR_TOTALBYTES_0), .Y(n3043) );
    zao2x4b U953 ( .A(DW1[31]), .B(n2652), .C(UP_DW5[4]), .D(n2291), .E(n2289), 
        .F(DW5[4]), .G(n2290), .H(NAKCNT996_3), .Y(NAKCNT1035_3) );
    zxo2b U954 ( .A(n2486), .B(n2485), .Y(NAKCNT996_3) );
    zao2x4b U955 ( .A(DW1[30]), .B(n2652), .C(UP_DW5[3]), .D(n2291), .E(n2289), 
        .F(DW5[3]), .G(NAKCNT996_2), .H(n2290), .Y(NAKCNT1035_2) );
    zxo2b U956 ( .A(UP_DW5[3]), .B(n2484), .Y(NAKCNT996_2) );
    zivb U957 ( .A(n2489), .Y(n2484) );
    zao2x4b U958 ( .A(DW1[29]), .B(n2652), .C(UP_DW5[2]), .D(n2291), .E(n2289), 
        .F(DW5[2]), .G(NAKCNT996_1), .H(n2290), .Y(NAKCNT1035_1) );
    znd2b U959 ( .A(n2489), .B(n2488), .Y(NAKCNT996_1) );
    zao2x4b U960 ( .A(DW1[28]), .B(n2652), .C(UP_DW5[1]), .D(n2291), .E(n2289), 
        .F(DW5[1]), .G(NAKCNT996_0), .H(n2290), .Y(NAKCNT1035_0) );
    zivb U961 ( .A(n3026), .Y(n3030) );
    zivb U962 ( .A(n3082), .Y(n3086) );
    zhadrb add_503_U1_1_1 ( .A(CPAGE_1), .B(CPAGE_0), .CO(add_503_carry_2), 
        .S(CPAGE1102_1) );
    zivb U963 ( .A(n3092), .Y(n3091) );
    zivb U964 ( .A(n2662), .Y(n3104) );
    zoai2x4b U965 ( .A(n2535), .B(n3159), .C(n2537), .D(n2538), .E(n2539), .F(
        n3161), .G(n2541), .H(n3163), .Y(CURQTDPTR1422_31) );
    zivb U966 ( .A(DW3[31]), .Y(n2535) );
    zivb U967 ( .A(DW4[31]), .Y(n2539) );
    zoai2x4b U968 ( .A(n2543), .B(n3158), .C(n3160), .D(n2544), .E(n2545), .F(
        n3162), .G(n2546), .H(n3164), .Y(CURQTDPTR1422_30) );
    zivb U969 ( .A(DW3[30]), .Y(n2543) );
    zivb U970 ( .A(DW4[30]), .Y(n2545) );
    zivb U971 ( .A(DW3[29]), .Y(n2547) );
    zivb U972 ( .A(DW4[29]), .Y(n2549) );
    zoai2x4b U973 ( .A(n2551), .B(n3159), .C(n3160), .D(n2552), .E(n2553), .F(
        n3161), .G(n2554), .H(n3163), .Y(CURQTDPTR1422_28) );
    zivb U974 ( .A(DW3[28]), .Y(n2551) );
    zivb U975 ( .A(DW4[28]), .Y(n2553) );
    zoai2x4b U976 ( .A(n2555), .B(n3158), .C(n2537), .D(n2556), .E(n2557), .F(
        n3162), .G(n2558), .H(n3164), .Y(CURQTDPTR1422_27) );
    zivb U977 ( .A(DW3[27]), .Y(n2555) );
    zivb U978 ( .A(DW4[27]), .Y(n2557) );
    zivb U979 ( .A(DW3[26]), .Y(n2559) );
    zivb U980 ( .A(DW4[26]), .Y(n2561) );
    zivb U981 ( .A(DW3[25]), .Y(n2563) );
    zivb U982 ( .A(DW4[25]), .Y(n2565) );
    zivb U983 ( .A(DW3[24]), .Y(n2567) );
    zivb U984 ( .A(DW4[24]), .Y(n2569) );
    zivb U985 ( .A(DW3[23]), .Y(n2571) );
    zivb U986 ( .A(DW4[23]), .Y(n2573) );
    zivb U987 ( .A(DW3[22]), .Y(n2575) );
    zivb U988 ( .A(DW4[22]), .Y(n2577) );
    zivb U989 ( .A(DW3[21]), .Y(n2579) );
    zivb U990 ( .A(DW4[21]), .Y(n2581) );
    zoai2x4b U991 ( .A(n2583), .B(n2536), .C(n3160), .D(n2584), .E(n2585), .F(
        n2540), .G(n2586), .H(n2542), .Y(CURQTDPTR1422_20) );
    zivb U992 ( .A(DW3[20]), .Y(n2583) );
    zivb U993 ( .A(DW4[20]), .Y(n2585) );
    zivb U994 ( .A(DW3[19]), .Y(n2587) );
    zivb U995 ( .A(DW4[19]), .Y(n2589) );
    zivb U996 ( .A(DW3[18]), .Y(n2591) );
    zivb U997 ( .A(DW4[18]), .Y(n2593) );
    zivb U998 ( .A(DW3[17]), .Y(n2595) );
    zivb U999 ( .A(DW4[17]), .Y(n2597) );
    zoai2x4b U1000 ( .A(n2599), .B(n3158), .C(n3160), .D(n2600), .E(n2601), 
        .F(n3161), .G(n2602), .H(n3163), .Y(CURQTDPTR1422_16) );
    zivb U1001 ( .A(DW3[16]), .Y(n2599) );
    zivb U1002 ( .A(DW4[16]), .Y(n2601) );
    zoai2x4b U1003 ( .A(n2603), .B(n3159), .C(n2537), .D(n2604), .E(n2605), 
        .F(n3162), .G(n2606), .H(n3164), .Y(CURQTDPTR1422_15) );
    zivb U1004 ( .A(DW3[15]), .Y(n2603) );
    zivb U1005 ( .A(DW4[15]), .Y(n2605) );
    zivb U1006 ( .A(DW3[14]), .Y(n2607) );
    zivb U1007 ( .A(DW4[14]), .Y(n2609) );
    zivb U1008 ( .A(DW3[13]), .Y(n2611) );
    zivb U1009 ( .A(DW4[13]), .Y(n2613) );
    zivb U1010 ( .A(DW3[12]), .Y(n2615) );
    zivb U1011 ( .A(DW4[12]), .Y(n2617) );
    zivb U1012 ( .A(DW3[11]), .Y(n2619) );
    zivb U1013 ( .A(DW4[11]), .Y(n2621) );
    zivb U1014 ( .A(DW5[11]), .Y(n2622) );
    zivb U1015 ( .A(DW3[10]), .Y(n2623) );
    zivb U1016 ( .A(DW4[10]), .Y(n2625) );
    zivb U1017 ( .A(DW5[10]), .Y(n2626) );
    zivb U1018 ( .A(DW3[9]), .Y(n2627) );
    zivb U1019 ( .A(DW4[9]), .Y(n2629) );
    zivb U1020 ( .A(DW5[9]), .Y(n2630) );
    zoai2x4b U1021 ( .A(n2631), .B(n2536), .C(n3160), .D(n2632), .E(n2633), 
        .F(n2540), .G(n2634), .H(n2542), .Y(CURQTDPTR1422_8) );
    zivb U1022 ( .A(DW3[8]), .Y(n2631) );
    zivb U1023 ( .A(DW4[8]), .Y(n2633) );
    zivb U1024 ( .A(DW5[8]), .Y(n2634) );
    zivb U1025 ( .A(DW3[7]), .Y(n2635) );
    zivb U1026 ( .A(DW4[7]), .Y(n2637) );
    zivb U1027 ( .A(DW5[7]), .Y(n2638) );
    zivb U1028 ( .A(DW3[6]), .Y(n2639) );
    zivb U1029 ( .A(DW4[6]), .Y(n2641) );
    zivb U1030 ( .A(DW5[6]), .Y(n2642) );
    zoai2x4b U1031 ( .A(n2643), .B(n2536), .C(n2537), .D(n2644), .E(n2645), 
        .F(n2540), .G(n2646), .H(n2542), .Y(CURQTDPTR1422_5) );
    zivb U1032 ( .A(DW3[5]), .Y(n2643) );
    zivb U1033 ( .A(n3088), .Y(n3090) );
    zivd U1034 ( .A(n3157), .Y(n2537) );
    zor2b U1035 ( .A(n2650), .B(n2534), .Y(n3157) );
    zivb U1036 ( .A(DW4[5]), .Y(n2645) );
    zivb U1037 ( .A(DW5[5]), .Y(n2646) );
    zivc U1038 ( .A(n3157), .Y(n3160) );
    zoai21b U1039 ( .A(n2505), .B(n2506), .C(n2320), .Y(PARSEQHEND_PRE) );
    zao21b U1040 ( .A(n2512), .B(QHSM[6]), .C(QHSM[9]), .Y(QEOT1815) );
    zivb U1041 ( .A(n2975), .Y(n2512) );
    zor2b U1042 ( .A(QCMDSTART), .B(n2514), .Y(n2975) );
    zmux21lb U1043 ( .A(n3019), .B(n2909), .S(n2320), .Y(SPLITXSTATE1256) );
    zmux21lb U1044 ( .A(n2502), .B(n3107), .S(n2320), .Y(ACTIVE_NXT) );
    zan2b U1045 ( .A(n2940), .B(n2941), .Y(n2761) );
    zivb U1046 ( .A(n2949), .Y(n2940) );
    zmux21lb U1047 ( .A(n2936), .B(n3100), .S(n2520), .Y(n2762) );
    zan3b U1048 ( .A(n2650), .B(n2534), .C(n2651), .Y(IMMEDRETRY1293) );
    zmux21lb U1049 ( .A(n3101), .B(n3052), .S(n2899), .Y(n2651) );
    zao33b U1050 ( .A(n2292), .B(n2501), .C(n2498), .D(n2297), .E(n2502), .F(
        n2503), .Y(QHSMNXT_1) );
    zivb U1051 ( .A(PCIEND), .Y(n2501) );
    zor2b U1052 ( .A(n3061), .B(n3060), .Y(n2503) );
    zivb U1053 ( .A(n3087), .Y(n3061) );
    zivb U1054 ( .A(DW4[0]), .Y(n3060) );
    zivb U1055 ( .A(QHSMNXT_1), .Y(n3089) );
    zivb U1056 ( .A(n2503), .Y(n2923) );
    znr3b U1057 ( .A(n2504), .B(ASYNC_EMPTY), .C(RECLAMATION), .Y(
        ASYNC_EMPTY1852) );
    zao21b U1058 ( .A(n3022), .B(n3023), .C(QRXERR), .Y(n2660) );
    zmux21lb U1059 ( .A(n2981), .B(n2898), .S(n2320), .Y(XACTERR1233) );
    zivb U1060 ( .A(n2660), .Y(n2900) );
    zivb U1061 ( .A(n2931), .Y(QHSMNXT_10) );
    znr2b U1062 ( .A(n2505), .B(n2513), .Y(CACHE_INVALID1602) );
    zan2b U1063 ( .A(n2533), .B(n2534), .Y(CACHE_MODIFY497) );
    zoai21b U1064 ( .A(LTINT_PCLK), .B(n2647), .C(n2648), .Y(QHIOCINT_T1889)
         );
    zivb U1065 ( .A(EHCI_MAC_EOT), .Y(n2514) );
    zoa211b U1066 ( .A(QHERRINT), .B(n2527), .C(n2528), .D(ERRINT_EN), .Y(
        QHERRINT2000) );
    znd2b U1067 ( .A(ERRINT), .B(LTINT_PCLK), .Y(n2528) );
    zoa211b U1068 ( .A(QHIOCINT), .B(n2529), .C(n2530), .D(USBINT_EN), .Y(
        QHIOCINT1926) );
    zoai21b U1069 ( .A(n2899), .B(n3063), .C(n3064), .Y(n2529) );
    zivc U1070 ( .A(n2521), .Y(n2899) );
    zivb U1071 ( .A(SPD), .Y(n3063) );
    znd2b U1072 ( .A(USBINT), .B(LTINT_PCLK), .Y(n2530) );
    zivb U1073 ( .A(n2529), .Y(n2648) );
    zivb U1074 ( .A(n2930), .Y(PHASENXT_resultwb) );
    znd2b U1075 ( .A(n2978), .B(n2498), .Y(n2930) );
    zoai21b U1076 ( .A(LTINT_PCLK), .B(n2531), .C(n2532), .Y(QHERRINT_T1963)
         );
    zivb U1077 ( .A(n2527), .Y(n2532) );
    zoai21b U1078 ( .A(n2656), .B(n2657), .C(n2658), .Y(DT881) );
    zivb U1079 ( .A(DW1[14]), .Y(n2950) );
    zivb U1080 ( .A(DW6[31]), .Y(n2657) );
    zmux21lb U1081 ( .A(n3103), .B(n3105), .S(UP_DW6[31]), .Y(n2658) );
    zivb U1082 ( .A(n2943), .Y(PING_PRESERVE) );
    zan2b U1083 ( .A(QHERRINT_T), .B(LTINT_PCLK), .Y(QHERRINT_S) );
    zan2b U1084 ( .A(LTINT_PCLK), .B(QHIOCINT_T), .Y(QHIOCINT_S) );
    zivb U1085 ( .A(n2504), .Y(HEADSEEN) );
    zivb U1086 ( .A(DW1[15]), .Y(n2967) );
    zivd U1087 ( .A(QH_PARSE_GO), .Y(n2534) );
    zao32b U1088 ( .A(n2496), .B(n2497), .C(n2498), .D(n2298), .E(TRAN_CMD
        [104]), .Y(QHSMNXT_7) );
    zivb U1089 ( .A(n2914), .Y(n2496) );
    zivb U1090 ( .A(QCMDSTART), .Y(n2497) );
    zivb U1091 ( .A(n3056), .Y(QHSMNXT_4) );
    znd2b U1092 ( .A(n3057), .B(n2498), .Y(n3056) );
    zao32b U1093 ( .A(n2499), .B(n2497), .C(n2498), .D(n2298), .E(n2500), .Y(
        QHSMNXT_5) );
    zivb U1094 ( .A(n2917), .Y(n2499) );
    zor2b U1095 ( .A(QHSM[8]), .B(QHSM[7]), .Y(n2508) );
    zivb U1096 ( .A(n2508), .Y(n3114) );
    zivb U1097 ( .A(n2659), .Y(QBUI_GO) );
    zan3b U1098 ( .A(UP_DW6[31]), .B(n2510), .C(n2511), .Y(TRAN_CMD[3]) );
    zivb U1099 ( .A(n2510), .Y(TRAN_CMD[7]) );
    zor2b U1100 ( .A(TRAN_CMD[9]), .B(n2522), .Y(n2510) );
    zan3b U1101 ( .A(n2522), .B(n2523), .C(n2511), .Y(TRAN_CMD[8]) );
    zivb U1102 ( .A(DW6[9]), .Y(n2522) );
    zivb U1103 ( .A(TRAN_CMD[9]), .Y(n2523) );
    zor2b U1104 ( .A(n2943), .B(n2939), .Y(n2511) );
    zivc U1105 ( .A(n2511), .Y(TRAN_CMD[5]) );
    zivb U1106 ( .A(DW1[27]), .Y(TRAN_CMD[11]) );
    zan2b U1107 ( .A(n2661), .B(MAXLEN[0]), .Y(TRAN_CMD[40]) );
    zan2b U1108 ( .A(n2661), .B(MAXLEN[1]), .Y(TRAN_CMD[41]) );
    zan2b U1109 ( .A(n2661), .B(MAXLEN[2]), .Y(TRAN_CMD[42]) );
    zan2b U1110 ( .A(n2661), .B(MAXLEN[3]), .Y(TRAN_CMD[43]) );
    zan2b U1111 ( .A(n2661), .B(MAXLEN[4]), .Y(TRAN_CMD[44]) );
    zan2b U1112 ( .A(n2661), .B(MAXLEN[5]), .Y(TRAN_CMD[45]) );
    zan2b U1113 ( .A(n2661), .B(MAXLEN[6]), .Y(TRAN_CMD[46]) );
    zan2b U1114 ( .A(n2661), .B(MAXLEN[7]), .Y(TRAN_CMD[47]) );
    zan2b U1115 ( .A(n2661), .B(MAXLEN[8]), .Y(TRAN_CMD[48]) );
    zan2b U1116 ( .A(n2661), .B(MAXLEN[9]), .Y(TRAN_CMD[49]) );
    zan2b U1117 ( .A(n2661), .B(MAXLEN[10]), .Y(TRAN_CMD[50]) );
    zivb U1118 ( .A(n2896), .Y(n3025) );
    zoai2x4b U1119 ( .A(n2326), .B(n2805), .C(n2806), .D(n2807), .E(n3169), 
        .F(n2809), .G(n2810), .H(n2811), .Y(TRAN_CMD[52]) );
    zivb U1120 ( .A(DW11[12]), .Y(n2811) );
    zoai2x4b U1121 ( .A(n2326), .B(n2812), .C(n3167), .D(n2813), .E(n2808), 
        .F(n2814), .G(n2810), .H(n2815), .Y(TRAN_CMD[53]) );
    zivb U1122 ( .A(DW11[13]), .Y(n2815) );
    zoai2x4b U1123 ( .A(n2326), .B(n2816), .C(n3166), .D(n2817), .E(n3168), 
        .F(n2818), .G(n2810), .H(n2819), .Y(TRAN_CMD[54]) );
    zivb U1124 ( .A(DW11[14]), .Y(n2819) );
    zoai2x4b U1125 ( .A(n2804), .B(n2820), .C(n2806), .D(n2821), .E(n3169), 
        .F(n2822), .G(n2810), .H(n2823), .Y(TRAN_CMD[55]) );
    zivb U1126 ( .A(DW11[15]), .Y(n2823) );
    zoai2x4b U1127 ( .A(n2326), .B(n2824), .C(n3167), .D(n2825), .E(n2808), 
        .F(n2826), .G(n2810), .H(n2827), .Y(TRAN_CMD[56]) );
    zivb U1128 ( .A(DW11[16]), .Y(n2827) );
    zoai2x4b U1129 ( .A(n2326), .B(n2828), .C(n2806), .D(n2829), .E(n3168), 
        .F(n2830), .G(n2810), .H(n2831), .Y(TRAN_CMD[57]) );
    zivb U1130 ( .A(DW11[17]), .Y(n2831) );
    zoai2x4b U1131 ( .A(n2804), .B(n2832), .C(n3166), .D(n2833), .E(n3169), 
        .F(n2834), .G(n2810), .H(n2835), .Y(TRAN_CMD[58]) );
    zivb U1132 ( .A(DW11[18]), .Y(n2835) );
    zoai2x4b U1133 ( .A(n2804), .B(n2836), .C(n3167), .D(n2837), .E(n2808), 
        .F(n2838), .G(n2810), .H(n2839), .Y(TRAN_CMD[59]) );
    zivb U1134 ( .A(DW11[19]), .Y(n2839) );
    zoai2x4b U1135 ( .A(n2804), .B(n2840), .C(n2806), .D(n2841), .E(n3168), 
        .F(n2842), .G(n2810), .H(n2843), .Y(TRAN_CMD[60]) );
    zivb U1136 ( .A(DW11[20]), .Y(n2843) );
    zoai2x4b U1137 ( .A(n2326), .B(n2844), .C(n3166), .D(n2845), .E(n3169), 
        .F(n2846), .G(n2810), .H(n2847), .Y(TRAN_CMD[61]) );
    zivb U1138 ( .A(DW11[21]), .Y(n2847) );
    zoai2x4b U1139 ( .A(n2326), .B(n2848), .C(n3166), .D(n2849), .E(n2808), 
        .F(n2850), .G(n2810), .H(n2851), .Y(TRAN_CMD[62]) );
    zivb U1140 ( .A(DW11[22]), .Y(n2851) );
    zoai2x4b U1141 ( .A(n2804), .B(n2852), .C(n3167), .D(n2853), .E(n3168), 
        .F(n2854), .G(n2810), .H(n2855), .Y(TRAN_CMD[63]) );
    zivb U1142 ( .A(DW11[23]), .Y(n2855) );
    zoai2x4b U1143 ( .A(n2326), .B(n2856), .C(n2806), .D(n2857), .E(n3169), 
        .F(n2858), .G(n2810), .H(n2859), .Y(TRAN_CMD[64]) );
    zivb U1144 ( .A(DW11[24]), .Y(n2859) );
    zoai2x4b U1145 ( .A(n2804), .B(n2860), .C(n3166), .D(n2861), .E(n2808), 
        .F(n2862), .G(n2810), .H(n2863), .Y(TRAN_CMD[65]) );
    zivb U1146 ( .A(DW11[25]), .Y(n2863) );
    zoai2x4b U1147 ( .A(n2804), .B(n2864), .C(n3167), .D(n2865), .E(n3168), 
        .F(n2866), .G(n2810), .H(n2867), .Y(TRAN_CMD[66]) );
    zivb U1148 ( .A(DW11[26]), .Y(n2867) );
    zoai2x4b U1149 ( .A(n2868), .B(n2326), .C(n2869), .D(n3166), .E(n2870), 
        .F(n2808), .G(n2810), .H(n2871), .Y(TRAN_CMD[67]) );
    zivb U1150 ( .A(DW11[27]), .Y(n2871) );
    zoai2x4b U1151 ( .A(n2804), .B(n2872), .C(n2806), .D(n2873), .E(n3169), 
        .F(n2874), .G(n2810), .H(n2875), .Y(TRAN_CMD[68]) );
    zivb U1152 ( .A(DW11[28]), .Y(n2875) );
    zoai2x4b U1153 ( .A(n2326), .B(n2876), .C(n3167), .D(n2877), .E(n2808), 
        .F(n2878), .G(n2810), .H(n2879), .Y(TRAN_CMD[69]) );
    zivb U1154 ( .A(DW11[29]), .Y(n2879) );
    zoai2x4b U1155 ( .A(n2804), .B(n2880), .C(n3166), .D(n2881), .E(n3168), 
        .F(n2882), .G(n2810), .H(n2883), .Y(TRAN_CMD[70]) );
    zivb U1156 ( .A(DW11[30]), .Y(n2883) );
    zoai2x4b U1157 ( .A(n2804), .B(n2884), .C(n2806), .D(n2885), .E(n3169), 
        .F(n2886), .G(n2810), .H(n2887), .Y(TRAN_CMD[71]) );
    zivf U1158 ( .A(n3152), .Y(n2810) );
    zao21b U1159 ( .A(CPAGE_0), .B(CPAGE_1), .C(n2328), .Y(n3152) );
    zivb U1160 ( .A(DW11[31]), .Y(n2887) );
    zan2b U1161 ( .A(DW8[12]), .B(n2902), .Y(n2802) );
    zan2b U1162 ( .A(DW8[13]), .B(n2902), .Y(n2800) );
    zan2b U1163 ( .A(DW8[14]), .B(n2902), .Y(n2798) );
    zan2b U1164 ( .A(DW8[15]), .B(n2902), .Y(n2796) );
    zan2b U1165 ( .A(DW8[16]), .B(n2902), .Y(n2794) );
    zan2b U1166 ( .A(DW8[17]), .B(n2902), .Y(n2792) );
    zan2b U1167 ( .A(DW8[18]), .B(n2902), .Y(n2790) );
    zan2b U1168 ( .A(DW8[19]), .B(n2902), .Y(n2788) );
    zan2b U1169 ( .A(DW8[20]), .B(n2902), .Y(n2786) );
    zan2b U1170 ( .A(DW8[21]), .B(n2902), .Y(n2784) );
    zan2b U1171 ( .A(DW8[22]), .B(n2902), .Y(n2782) );
    zan2b U1172 ( .A(DW8[23]), .B(n2902), .Y(n2780) );
    zan2b U1173 ( .A(DW8[24]), .B(n2902), .Y(n2778) );
    zan2b U1174 ( .A(DW8[25]), .B(n2902), .Y(n2776) );
    zan2b U1175 ( .A(DW8[26]), .B(n2902), .Y(n2774) );
    zan2b U1176 ( .A(n2902), .B(DW8[27]), .Y(n2772) );
    zan2b U1177 ( .A(DW8[28]), .B(n2902), .Y(n2770) );
    zan2b U1178 ( .A(DW8[29]), .B(n2902), .Y(n2768) );
    zan2b U1179 ( .A(DW8[30]), .B(n2902), .Y(n2766) );
    zivf U1180 ( .A(n3165), .Y(n2763) );
    zan2b U1181 ( .A(DW8[31]), .B(n2902), .Y(n2764) );
    zivf U1182 ( .A(n3167), .Y(n2902) );
    zivf U1183 ( .A(n3020), .Y(n3109) );
    zivf U1184 ( .A(n3168), .Y(n3110) );
    zor2b U1185 ( .A(UP_DW6[8]), .B(n2524), .Y(TRAN_CMD[104]) );
    zivb U1186 ( .A(n3021), .Y(n2524) );
    zor2b U1187 ( .A(n2515), .B(n2910), .Y(n3021) );
    zivb U1188 ( .A(TRAN_CMD[6]), .Y(n2515) );
    zivb U1189 ( .A(TRAN_CMD[104]), .Y(n2500) );
    zao22b U1190 ( .A(DW11[0]), .B(n3176), .C(DW6[0]), .D(n3127), .Y(n2666) );
    zao2x4b U1191 ( .A(DW5[0]), .B(n3128), .C(DW8[0]), .D(n3129), .E(DW9[0]), 
        .F(n3130), .G(DW10[0]), .H(n3131), .Y(n2667) );
    zao22b U1192 ( .A(DW11[1]), .B(n3126), .C(DW6[1]), .D(n3178), .Y(n2669) );
    zao2x4b U1193 ( .A(DW5[1]), .B(n3128), .C(DW8[1]), .D(n3129), .E(DW9[1]), 
        .F(n3130), .G(DW10[1]), .H(n3131), .Y(n2670) );
    zao22b U1194 ( .A(DW11[2]), .B(n3176), .C(DW6[2]), .D(n3127), .Y(n2672) );
    zao2x4b U1195 ( .A(DW5[2]), .B(n3128), .C(DW8[2]), .D(n3129), .E(DW9[2]), 
        .F(n3130), .G(DW10[2]), .H(n3131), .Y(n2673) );
    zao22b U1196 ( .A(DW11[3]), .B(n3126), .C(DW6[3]), .D(n3177), .Y(n2675) );
    zao2x4b U1197 ( .A(DW5[3]), .B(n3128), .C(DW8[3]), .D(n3129), .E(DW9[3]), 
        .F(n3130), .G(DW10[3]), .H(n3131), .Y(n2676) );
    zao22b U1198 ( .A(DW11[4]), .B(n3176), .C(DW6[4]), .D(n3177), .Y(n2678) );
    zao2x4b U1199 ( .A(DW5[4]), .B(n3128), .C(DW8[4]), .D(n3129), .E(DW9[4]), 
        .F(n3130), .G(DW10[4]), .H(n3131), .Y(n2679) );
    zao22b U1200 ( .A(DW11[5]), .B(n3126), .C(DW6[5]), .D(n3127), .Y(n2681) );
    zao2x4b U1201 ( .A(DW5[5]), .B(n3128), .C(DW8[5]), .D(n3129), .E(DW9[5]), 
        .F(n3130), .G(DW10[5]), .H(n3131), .Y(n2682) );
    zao22b U1202 ( .A(DW11[6]), .B(n3176), .C(DW6[6]), .D(n3178), .Y(n2684) );
    zao2x4b U1203 ( .A(DW5[6]), .B(n3128), .C(DW8[6]), .D(n3129), .E(DW9[6]), 
        .F(n3130), .G(DW10[6]), .H(n3131), .Y(n2685) );
    zao22b U1204 ( .A(DW11[7]), .B(n3126), .C(DW6[7]), .D(n3177), .Y(n2687) );
    zao2x4b U1205 ( .A(DW5[7]), .B(n3128), .C(DW8[7]), .D(n3129), .E(DW9[7]), 
        .F(n3130), .G(DW10[7]), .H(n3131), .Y(n2688) );
    zao22b U1206 ( .A(DW11[8]), .B(n3176), .C(TRAN_CMD[9]), .D(n3127), .Y(
        n2690) );
    zbfd U1207 ( .A(DW6[8]), .Y(TRAN_CMD[9]) );
    zao2x4b U1208 ( .A(DW5[8]), .B(n3128), .C(DW8[8]), .D(n3129), .E(DW9[8]), 
        .F(n3130), .G(DW10[8]), .H(n3131), .Y(n2691) );
    zao22b U1209 ( .A(n3126), .B(DW11[9]), .C(DW6[9]), .D(n3178), .Y(n2693) );
    zao2x4b U1210 ( .A(n3128), .B(DW5[9]), .C(n3129), .D(DW8[9]), .E(n3130), 
        .F(DW9[9]), .G(n3131), .H(DW10[9]), .Y(n2694) );
    zao22b U1211 ( .A(DW11[10]), .B(n3176), .C(DW6[10]), .D(n3177), .Y(n2696)
         );
    zao2x4b U1212 ( .A(DW5[10]), .B(n3128), .C(DW8[10]), .D(n3129), .E(DW9[10]
        ), .F(n3130), .G(DW10[10]), .H(n3131), .Y(n2697) );
    zao22b U1213 ( .A(DW11[11]), .B(n3126), .C(DW6[11]), .D(n3127), .Y(n2699)
         );
    zao2x4b U1214 ( .A(DW5[11]), .B(n3128), .C(DW8[11]), .D(n3129), .E(DW9[11]
        ), .F(n3130), .G(DW10[11]), .H(n3131), .Y(n2700) );
    zivc U1215 ( .A(n3079), .Y(n3128) );
    zivc U1216 ( .A(n3078), .Y(n3129) );
    zivc U1217 ( .A(n3183), .Y(n3130) );
    zivc U1218 ( .A(n3186), .Y(n3131) );
    zao22b U1219 ( .A(n3126), .B(DW11[12]), .C(DW6[12]), .D(n3178), .Y(n2702)
         );
    zoai2x4b U1220 ( .A(n3180), .B(n2618), .C(n2805), .D(n3078), .E(n2807), 
        .F(n3077), .G(n2809), .H(n3076), .Y(n2703) );
    zivb U1221 ( .A(DW5[12]), .Y(n2618) );
    zivb U1222 ( .A(DW8[12]), .Y(n2805) );
    zivb U1223 ( .A(DW9[12]), .Y(n2807) );
    zivb U1224 ( .A(DW10[12]), .Y(n2809) );
    zao22b U1225 ( .A(n3176), .B(DW11[13]), .C(DW6[13]), .D(n3177), .Y(n2705)
         );
    zoai2x4b U1226 ( .A(n3179), .B(n2614), .C(n2812), .D(n3182), .E(n2813), 
        .F(n3184), .G(n2814), .H(n3186), .Y(n2706) );
    zivb U1227 ( .A(DW5[13]), .Y(n2614) );
    zivb U1228 ( .A(DW8[13]), .Y(n2812) );
    zivb U1229 ( .A(DW9[13]), .Y(n2813) );
    zivb U1230 ( .A(DW10[13]), .Y(n2814) );
    zao22b U1231 ( .A(n3126), .B(DW11[14]), .C(DW6[14]), .D(n3127), .Y(n2708)
         );
    zoai2x4b U1232 ( .A(n3079), .B(n2610), .C(n2816), .D(n3181), .E(n2817), 
        .F(n3183), .G(n2818), .H(n3185), .Y(n2709) );
    zivb U1233 ( .A(DW5[14]), .Y(n2610) );
    zivb U1234 ( .A(DW8[14]), .Y(n2816) );
    zivb U1235 ( .A(DW9[14]), .Y(n2817) );
    zivb U1236 ( .A(DW10[14]), .Y(n2818) );
    zao22b U1237 ( .A(n3176), .B(DW11[15]), .C(DW6[15]), .D(n3178), .Y(n2711)
         );
    zoai2x4b U1238 ( .A(n3180), .B(n2606), .C(n2820), .D(n3182), .E(n2821), 
        .F(n3077), .G(n2822), .H(n3076), .Y(n2712) );
    zivb U1239 ( .A(DW5[15]), .Y(n2606) );
    zivb U1240 ( .A(DW8[15]), .Y(n2820) );
    zivb U1241 ( .A(DW9[15]), .Y(n2821) );
    zivb U1242 ( .A(DW10[15]), .Y(n2822) );
    zao22b U1243 ( .A(n3126), .B(DW11[16]), .C(DW6[16]), .D(n3177), .Y(n2714)
         );
    zoai2x4b U1244 ( .A(n3179), .B(n2602), .C(n2824), .D(n3181), .E(n2825), 
        .F(n3184), .G(n2826), .H(n3185), .Y(n2715) );
    zivb U1245 ( .A(DW5[16]), .Y(n2602) );
    zivb U1246 ( .A(DW8[16]), .Y(n2824) );
    zivb U1247 ( .A(DW9[16]), .Y(n2825) );
    zivb U1248 ( .A(DW10[16]), .Y(n2826) );
    zao22b U1249 ( .A(n3176), .B(DW11[17]), .C(DW6[17]), .D(n3127), .Y(n2717)
         );
    zoai2x4b U1250 ( .A(n3079), .B(n2598), .C(n2828), .D(n3078), .E(n2829), 
        .F(n3183), .G(n2830), .H(n3186), .Y(n2718) );
    zivb U1251 ( .A(DW5[17]), .Y(n2598) );
    zivb U1252 ( .A(DW8[17]), .Y(n2828) );
    zivb U1253 ( .A(DW9[17]), .Y(n2829) );
    zivb U1254 ( .A(DW10[17]), .Y(n2830) );
    zao22b U1255 ( .A(n3126), .B(DW11[18]), .C(DW6[18]), .D(n3178), .Y(n2720)
         );
    zoai2x4b U1256 ( .A(n3180), .B(n2594), .C(n2832), .D(n3182), .E(n2833), 
        .F(n3077), .G(n2834), .H(n3076), .Y(n2721) );
    zivb U1257 ( .A(DW5[18]), .Y(n2594) );
    zivb U1258 ( .A(DW8[18]), .Y(n2832) );
    zivb U1259 ( .A(DW9[18]), .Y(n2833) );
    zivb U1260 ( .A(DW10[18]), .Y(n2834) );
    zao22b U1261 ( .A(n3176), .B(DW11[19]), .C(DW6[19]), .D(n3177), .Y(n2723)
         );
    zoai2x4b U1262 ( .A(n3179), .B(n2590), .C(n2836), .D(n3181), .E(n2837), 
        .F(n3184), .G(n2838), .H(n3186), .Y(n2724) );
    zivb U1263 ( .A(DW5[19]), .Y(n2590) );
    zivb U1264 ( .A(DW8[19]), .Y(n2836) );
    zivb U1265 ( .A(DW9[19]), .Y(n2837) );
    zivb U1266 ( .A(DW10[19]), .Y(n2838) );
    zao22b U1267 ( .A(n3126), .B(DW11[20]), .C(DW6[20]), .D(n3178), .Y(n2726)
         );
    zoai2x4b U1268 ( .A(n3079), .B(n2586), .C(n2840), .D(n3078), .E(n2841), 
        .F(n3183), .G(n2842), .H(n3185), .Y(n2727) );
    zivb U1269 ( .A(DW5[20]), .Y(n2586) );
    zivb U1270 ( .A(DW8[20]), .Y(n2840) );
    zivb U1271 ( .A(DW9[20]), .Y(n2841) );
    zivb U1272 ( .A(DW10[20]), .Y(n2842) );
    zao22b U1273 ( .A(n3176), .B(DW11[21]), .C(DW6[21]), .D(n3177), .Y(n2729)
         );
    zoai2x4b U1274 ( .A(n3180), .B(n2582), .C(n2844), .D(n3182), .E(n2845), 
        .F(n3077), .G(n2846), .H(n3076), .Y(n2730) );
    zivb U1275 ( .A(DW5[21]), .Y(n2582) );
    zivb U1276 ( .A(DW8[21]), .Y(n2844) );
    zivb U1277 ( .A(DW9[21]), .Y(n2845) );
    zivb U1278 ( .A(DW10[21]), .Y(n2846) );
    zao22b U1279 ( .A(n3126), .B(DW11[22]), .C(DW6[22]), .D(n3127), .Y(n2732)
         );
    zoai2x4b U1280 ( .A(n3179), .B(n2578), .C(n2848), .D(n3181), .E(n2849), 
        .F(n3184), .G(n2850), .H(n3186), .Y(n2733) );
    zivb U1281 ( .A(DW5[22]), .Y(n2578) );
    zivb U1282 ( .A(DW8[22]), .Y(n2848) );
    zivb U1283 ( .A(DW9[22]), .Y(n2849) );
    zivb U1284 ( .A(DW10[22]), .Y(n2850) );
    zao22b U1285 ( .A(n3176), .B(DW11[23]), .C(DW6[23]), .D(n3178), .Y(n2735)
         );
    zoai2x4b U1286 ( .A(n3079), .B(n2574), .C(n2852), .D(n3078), .E(n2853), 
        .F(n3183), .G(n2854), .H(n3185), .Y(n2736) );
    zivb U1287 ( .A(DW5[23]), .Y(n2574) );
    zivb U1288 ( .A(DW8[23]), .Y(n2852) );
    zivb U1289 ( .A(DW9[23]), .Y(n2853) );
    zivb U1290 ( .A(DW10[23]), .Y(n2854) );
    zao22b U1291 ( .A(n3126), .B(DW11[24]), .C(DW6[24]), .D(n3177), .Y(n2738)
         );
    zoai2x4b U1292 ( .A(n3180), .B(n2570), .C(n2856), .D(n3182), .E(n2857), 
        .F(n3077), .G(n2858), .H(n3076), .Y(n2739) );
    zivb U1293 ( .A(DW5[24]), .Y(n2570) );
    zivb U1294 ( .A(DW8[24]), .Y(n2856) );
    zivb U1295 ( .A(DW9[24]), .Y(n2857) );
    zivb U1296 ( .A(DW10[24]), .Y(n2858) );
    zao22b U1297 ( .A(n3176), .B(DW11[25]), .C(DW6[25]), .D(n3127), .Y(n2741)
         );
    zoai2x4b U1298 ( .A(n3179), .B(n2566), .C(n2860), .D(n3181), .E(n2861), 
        .F(n3184), .G(n2862), .H(n3186), .Y(n2742) );
    zivb U1299 ( .A(DW5[25]), .Y(n2566) );
    zivb U1300 ( .A(DW8[25]), .Y(n2860) );
    zivb U1301 ( .A(DW9[25]), .Y(n2861) );
    zivb U1302 ( .A(DW10[25]), .Y(n2862) );
    zao22b U1303 ( .A(n3126), .B(DW11[26]), .C(DW6[26]), .D(n3178), .Y(n2744)
         );
    zoai2x4b U1304 ( .A(n3079), .B(n2562), .C(n2864), .D(n3078), .E(n2865), 
        .F(n3183), .G(n2866), .H(n3185), .Y(n2745) );
    zivb U1305 ( .A(DW5[26]), .Y(n2562) );
    zivb U1306 ( .A(DW8[26]), .Y(n2864) );
    zivb U1307 ( .A(DW9[26]), .Y(n2865) );
    zivb U1308 ( .A(DW10[26]), .Y(n2866) );
    zao22b U1309 ( .A(n3176), .B(DW11[27]), .C(DW6[27]), .D(n3177), .Y(n2747)
         );
    zoai2x4b U1310 ( .A(n3180), .B(n2558), .C(n2868), .D(n3182), .E(n2869), 
        .F(n3077), .G(n2870), .H(n3076), .Y(n2748) );
    zivb U1311 ( .A(DW5[27]), .Y(n2558) );
    zivb U1312 ( .A(DW8[27]), .Y(n2868) );
    zivb U1313 ( .A(DW9[27]), .Y(n2869) );
    zivb U1314 ( .A(DW10[27]), .Y(n2870) );
    zao22b U1315 ( .A(n3126), .B(DW11[28]), .C(DW6[28]), .D(n3127), .Y(n2750)
         );
    zoai2x4b U1316 ( .A(n3179), .B(n2554), .C(n2872), .D(n3181), .E(n2873), 
        .F(n3184), .G(n2874), .H(n3186), .Y(n2751) );
    zivb U1317 ( .A(DW5[28]), .Y(n2554) );
    zivb U1318 ( .A(DW8[28]), .Y(n2872) );
    zivb U1319 ( .A(DW9[28]), .Y(n2873) );
    zivb U1320 ( .A(DW10[28]), .Y(n2874) );
    zao22b U1321 ( .A(n3176), .B(DW11[29]), .C(DW6[29]), .D(n3178), .Y(n2753)
         );
    zoai2x4b U1322 ( .A(n3079), .B(n2550), .C(n2876), .D(n3078), .E(n2877), 
        .F(n3183), .G(n2878), .H(n3185), .Y(n2754) );
    zivb U1323 ( .A(DW5[29]), .Y(n2550) );
    zivb U1324 ( .A(DW8[29]), .Y(n2876) );
    zivb U1325 ( .A(DW9[29]), .Y(n2877) );
    zivb U1326 ( .A(DW10[29]), .Y(n2878) );
    zivd U1327 ( .A(n3068), .Y(n3124) );
    zao22b U1328 ( .A(n3126), .B(DW11[30]), .C(DW6[30]), .D(n3127), .Y(n2756)
         );
    zivd U1329 ( .A(n3075), .Y(n3126) );
    zoai2x4b U1330 ( .A(n3180), .B(n2546), .C(n2880), .D(n3182), .E(n2881), 
        .F(n3077), .G(n2882), .H(n3076), .Y(n2757) );
    zivb U1331 ( .A(DW5[30]), .Y(n2546) );
    zivb U1332 ( .A(DW8[30]), .Y(n2880) );
    zivb U1333 ( .A(DW9[30]), .Y(n2881) );
    zivb U1334 ( .A(DW10[30]), .Y(n2882) );
    zivd U1335 ( .A(n3068), .Y(n3173) );
    zao22b U1336 ( .A(n3176), .B(DW11[31]), .C(DW6[31]), .D(n3178), .Y(n2759)
         );
    zivd U1337 ( .A(n3075), .Y(n3176) );
    zoai2x4b U1338 ( .A(n3179), .B(n2541), .C(n2884), .D(n3181), .E(n2885), 
        .F(n3184), .G(n2886), .H(n3185), .Y(n2760) );
    zivb U1339 ( .A(DW5[31]), .Y(n2541) );
    zivb U1340 ( .A(DW8[31]), .Y(n2884) );
    zivb U1341 ( .A(DW9[31]), .Y(n2885) );
    zivb U1342 ( .A(DW10[31]), .Y(n2886) );
    zmux21hb U1343 ( .A(UP_DW3[5]), .B(CACHE_ADDR[0]), .S(QHSM[12]), .Y(
        QHCIADR[5]) );
    zmux21hb U1344 ( .A(UP_DW3[6]), .B(CACHE_ADDR[1]), .S(QHSM[12]), .Y(
        QHCIADR[6]) );
    zmux21hb U1345 ( .A(UP_DW3[7]), .B(CACHE_ADDR[2]), .S(QHDWNUM[3]), .Y(
        QHCIADR[7]) );
    zmux21hb U1346 ( .A(UP_DW3[8]), .B(CACHE_ADDR[3]), .S(QHSM[12]), .Y(
        QHCIADR[8]) );
    zmux21hb U1347 ( .A(UP_DW3[9]), .B(CACHE_ADDR[4]), .S(n2358), .Y(QHCIADR
        [9]) );
    zmux21hb U1348 ( .A(UP_DW3[10]), .B(CACHE_ADDR[5]), .S(QHDWNUM[3]), .Y(
        QHCIADR[10]) );
    zmux21hb U1349 ( .A(UP_DW3[11]), .B(CACHE_ADDR[6]), .S(QHSM[12]), .Y(
        QHCIADR[11]) );
    zmux21hb U1350 ( .A(UP_DW3[12]), .B(CACHE_ADDR[7]), .S(QHDWNUM[3]), .Y(
        QHCIADR[12]) );
    zmux21hb U1351 ( .A(UP_DW3[13]), .B(CACHE_ADDR[8]), .S(QHSM[12]), .Y(
        QHCIADR[13]) );
    zmux21hb U1352 ( .A(UP_DW3[14]), .B(CACHE_ADDR[9]), .S(QHSM[12]), .Y(
        QHCIADR[14]) );
    zmux21hb U1353 ( .A(UP_DW3[15]), .B(CACHE_ADDR[10]), .S(QHDWNUM[3]), .Y(
        QHCIADR[15]) );
    zmux21hb U1354 ( .A(UP_DW3[16]), .B(CACHE_ADDR[11]), .S(QHDWNUM[3]), .Y(
        QHCIADR[16]) );
    zmux21hb U1355 ( .A(UP_DW3[17]), .B(CACHE_ADDR[12]), .S(QHDWNUM[3]), .Y(
        QHCIADR[17]) );
    zmux21hb U1356 ( .A(UP_DW3[18]), .B(CACHE_ADDR[13]), .S(QHDWNUM[3]), .Y(
        QHCIADR[18]) );
    zmux21hb U1357 ( .A(UP_DW3[19]), .B(CACHE_ADDR[14]), .S(QHCIADR[2]), .Y(
        QHCIADR[19]) );
    zmux21hb U1358 ( .A(UP_DW3[20]), .B(CACHE_ADDR[15]), .S(QHSM[12]), .Y(
        QHCIADR[20]) );
    zmux21hb U1359 ( .A(UP_DW3[21]), .B(CACHE_ADDR[16]), .S(QHSM[12]), .Y(
        QHCIADR[21]) );
    zmux21hb U1360 ( .A(UP_DW3[22]), .B(CACHE_ADDR[17]), .S(QHDWNUM[3]), .Y(
        QHCIADR[22]) );
    zmux21hb U1361 ( .A(UP_DW3[23]), .B(CACHE_ADDR[18]), .S(QHDWNUM[3]), .Y(
        QHCIADR[23]) );
    zmux21hb U1362 ( .A(UP_DW3[24]), .B(CACHE_ADDR[19]), .S(QHCIADR[2]), .Y(
        QHCIADR[24]) );
    zmux21hb U1363 ( .A(UP_DW3[25]), .B(CACHE_ADDR[20]), .S(QHDWNUM[3]), .Y(
        QHCIADR[25]) );
    zmux21hb U1364 ( .A(UP_DW3[26]), .B(CACHE_ADDR[21]), .S(QHCIADR[2]), .Y(
        QHCIADR[26]) );
    zmux21hb U1365 ( .A(UP_DW3[27]), .B(CACHE_ADDR[22]), .S(QHSM[12]), .Y(
        QHCIADR[27]) );
    zmux21hb U1366 ( .A(UP_DW3[28]), .B(CACHE_ADDR[23]), .S(QHDWNUM[3]), .Y(
        QHCIADR[28]) );
    zmux21hb U1367 ( .A(UP_DW3[29]), .B(CACHE_ADDR[24]), .S(QHDWNUM[3]), .Y(
        QHCIADR[29]) );
    zmux21hb U1368 ( .A(UP_DW3[30]), .B(CACHE_ADDR[25]), .S(QHDWNUM[3]), .Y(
        QHCIADR[30]) );
    zmux21hb U1369 ( .A(UP_DW3[31]), .B(CACHE_ADDR[26]), .S(QHDWNUM[3]), .Y(
        QHCIADR[31]) );
    zor2b U1370 ( .A(QHSM[1]), .B(QHCIMWR), .Y(QHCIREQ) );
    zor2b U1371 ( .A(QHSM[2]), .B(QHSM[11]), .Y(CACHEPHASE) );
    zmux21lb U1372 ( .A(n2910), .B(n3019), .S(n2525), .Y(UP_DW6[1]) );
    zivb U1373 ( .A(DW6[1]), .Y(n3019) );
    zan2b U1374 ( .A(DW6[2]), .B(n2525), .Y(UP_DW6[2]) );
    zmux21lb U1375 ( .A(n2901), .B(n2981), .S(n2525), .Y(UP_DW6[3]) );
    zivb U1376 ( .A(DW6[3]), .Y(n2981) );
    zao21b U1377 ( .A(BABBLE), .B(n2526), .C(DW6[4]), .Y(UP_DW6[4]) );
    zan2b U1378 ( .A(DW6[5]), .B(n3170), .Y(UP_DW6[5]) );
    zmux21lb U1379 ( .A(n3095), .B(n2982), .S(n2525), .Y(UP_DW6[6]) );
    zivb U1380 ( .A(DW6[6]), .Y(n2982) );
    zmux21lb U1381 ( .A(n2959), .B(n2502), .S(n3170), .Y(UP_DW6[7]) );
    zivb U1382 ( .A(DW6[7]), .Y(n2502) );
    zbfd U1383 ( .A(DW6[8]), .Y(UP_DW6[8]) );
    zmux21lb U1384 ( .A(n3045), .B(n3018), .S(n3170), .Y(UP_DW6[10]) );
    zivb U1385 ( .A(DW6[10]), .Y(n3018) );
    zmux21lb U1386 ( .A(n2490), .B(n3017), .S(n2525), .Y(UP_DW6[11]) );
    zivb U1387 ( .A(DW6[11]), .Y(n3017) );
    zmux21lb U1388 ( .A(n3016), .B(n3015), .S(n3170), .Y(UP_DW6[12]) );
    zivb U1389 ( .A(DW6[12]), .Y(n3015) );
    zmux21lb U1390 ( .A(n3014), .B(n3013), .S(n2525), .Y(UP_DW6[13]) );
    zivb U1391 ( .A(DW6[13]), .Y(n3013) );
    zmux21lb U1392 ( .A(n3012), .B(n3011), .S(n3170), .Y(UP_DW6[14]) );
    zivb U1393 ( .A(DW6[14]), .Y(n3011) );
    zmux21lb U1394 ( .A(n3010), .B(n3009), .S(n2525), .Y(UP_DW6[16]) );
    zivb U1395 ( .A(DW6[16]), .Y(n3009) );
    zmux21lb U1396 ( .A(n3008), .B(n3007), .S(n3170), .Y(UP_DW6[17]) );
    zivb U1397 ( .A(DW6[17]), .Y(n3007) );
    zmux21lb U1398 ( .A(n3006), .B(n3005), .S(n2525), .Y(UP_DW6[18]) );
    zivb U1399 ( .A(DW6[18]), .Y(n3005) );
    zmux21lb U1400 ( .A(n3004), .B(n3003), .S(n3170), .Y(UP_DW6[19]) );
    zivb U1401 ( .A(DW6[19]), .Y(n3003) );
    zmux21lb U1402 ( .A(n3002), .B(n3001), .S(n2525), .Y(UP_DW6[20]) );
    zivb U1403 ( .A(DW6[20]), .Y(n3001) );
    zmux21lb U1404 ( .A(n3000), .B(n2999), .S(n3170), .Y(UP_DW6[21]) );
    zivb U1405 ( .A(DW6[21]), .Y(n2999) );
    zmux21lb U1406 ( .A(n2998), .B(n2997), .S(n2525), .Y(UP_DW6[22]) );
    zivb U1407 ( .A(DW6[22]), .Y(n2997) );
    zmux21lb U1408 ( .A(n2996), .B(n2995), .S(n3170), .Y(UP_DW6[23]) );
    zivb U1409 ( .A(DW6[23]), .Y(n2995) );
    zmux21lb U1410 ( .A(n2994), .B(n2993), .S(n2525), .Y(UP_DW6[24]) );
    zivb U1411 ( .A(DW6[24]), .Y(n2993) );
    zmux21lb U1412 ( .A(n2992), .B(n2991), .S(n3170), .Y(UP_DW6[25]) );
    zivb U1413 ( .A(DW6[25]), .Y(n2991) );
    zmux21lb U1414 ( .A(n2990), .B(n2989), .S(n2525), .Y(UP_DW6[26]) );
    zivb U1415 ( .A(DW6[26]), .Y(n2989) );
    zmux21lb U1416 ( .A(n2429), .B(n2988), .S(n3170), .Y(UP_DW6[27]) );
    zivb U1417 ( .A(DW6[27]), .Y(n2988) );
    zmux21lb U1418 ( .A(n2428), .B(n2987), .S(n2525), .Y(UP_DW6[28]) );
    zivb U1419 ( .A(DW6[28]), .Y(n2987) );
    zmux21lb U1420 ( .A(n2986), .B(n2985), .S(n3170), .Y(UP_DW6[29]) );
    zivb U1421 ( .A(DW6[29]), .Y(n2985) );
    zmux21lb U1422 ( .A(n2984), .B(n2983), .S(n3170), .Y(UP_DW6[30]) );
    zivb U1423 ( .A(DW6[30]), .Y(n2983) );
    zivd U1424 ( .A(n2526), .Y(n3170) );
    zor2b U1425 ( .A(UP_LDW7), .B(QHSM[11]), .Y(n2526) );
    zivd U1426 ( .A(n2526), .Y(n2525) );
    znd2b U1427 ( .A(n3137), .B(n2498), .Y(n2517) );
    zivb U1428 ( .A(PHASENXT_idle), .Y(n2505) );
    zivb U1429 ( .A(n2969), .Y(n2491) );
    zor2b U1430 ( .A(n2929), .B(n3156), .Y(n2519) );
    zivb U1431 ( .A(n3101), .Y(n3156) );
    zivb U1432 ( .A(n2517), .Y(QHSMNXT_12) );
    zivb U1433 ( .A(n2518), .Y(QHSMNXT_13) );
    zivb U1434 ( .A(QHSM[3]), .Y(n3049) );
    zivc U1435 ( .A(QHSM[0]), .Y(n2650) );
    zdffqrb TOTALBYTES_reg_14 ( .CK(PCICLK), .D(TOTALBYTES640_14), .R(TRST_), 
        .Q(TOTALBYTES_14) );
    zivb U1436 ( .A(TOTALBYTES_14), .Y(n2984) );
    zdffqrb TOTALBYTES_reg_13 ( .CK(PCICLK), .D(TOTALBYTES640_13), .R(TRST_), 
        .Q(TOTALBYTES_13) );
    zivb U1437 ( .A(TOTALBYTES_13), .Y(n2986) );
    zdffqrb TOTALBYTES_reg_10 ( .CK(PCICLK), .D(TOTALBYTES640_10), .R(TRST_), 
        .Q(TOTALBYTES_10) );
    zivb U1438 ( .A(TOTALBYTES_10), .Y(n2990) );
    zdffqrb TOTALBYTES_reg_1 ( .CK(PCICLK), .D(TOTALBYTES640_1), .R(TRST_), 
        .Q(TOTALBYTES_1) );
    zivb U1439 ( .A(TOTALBYTES_1), .Y(n3008) );
    zdffqrb TOTALBYTES_reg_0 ( .CK(PCICLK), .D(TOTALBYTES640_0), .R(TRST_), 
        .Q(TOTALBYTES_0) );
    zivb U1440 ( .A(TOTALBYTES_0), .Y(n3010) );
    zdffrb NAKCNT_reg_3 ( .CK(PCICLK), .D(NAKCNT1035_3), .R(TRST_), .Q(UP_DW5
        [4]), .QN(n2486) );
    zdffqrb NAKCNT_reg_2 ( .CK(PCICLK), .D(NAKCNT1035_2), .R(TRST_), .Q(UP_DW5
        [3]) );
    zivb U1441 ( .A(UP_DW5[3]), .Y(n2483) );
    zdffqrb NAKCNT_reg_1 ( .CK(PCICLK), .D(NAKCNT1035_1), .R(TRST_), .Q(UP_DW5
        [2]) );
    zivb U1442 ( .A(UP_DW5[2]), .Y(n2487) );
    zdffqrb NAKCNT_reg_0 ( .CK(PCICLK), .D(NAKCNT1035_0), .R(TRST_), .Q(UP_DW5
        [1]) );
    zivb U1443 ( .A(UP_DW5[1]), .Y(NAKCNT996_0) );
    zivb U1444 ( .A(CPAGE_1), .Y(n3014) );
    zdffb CURQTDPTR_reg_31 ( .CK(PCICLK), .D(CURQTDPTR1422_31), .Q(UP_DW3[31]), 
        .QN(n2538) );
    zdffb CURQTDPTR_reg_30 ( .CK(PCICLK), .D(CURQTDPTR1422_30), .Q(UP_DW3[30]), 
        .QN(n2544) );
    zdffb CURQTDPTR_reg_29 ( .CK(PCICLK), .D(CURQTDPTR1422_29), .Q(UP_DW3[29]), 
        .QN(n2548) );
    zdffb CURQTDPTR_reg_28 ( .CK(PCICLK), .D(CURQTDPTR1422_28), .Q(UP_DW3[28]), 
        .QN(n2552) );
    zdffb CURQTDPTR_reg_27 ( .CK(PCICLK), .D(CURQTDPTR1422_27), .Q(UP_DW3[27]), 
        .QN(n2556) );
    zdffb CURQTDPTR_reg_26 ( .CK(PCICLK), .D(CURQTDPTR1422_26), .Q(UP_DW3[26]), 
        .QN(n2560) );
    zdffb CURQTDPTR_reg_25 ( .CK(PCICLK), .D(CURQTDPTR1422_25), .Q(UP_DW3[25]), 
        .QN(n2564) );
    zdffb CURQTDPTR_reg_24 ( .CK(PCICLK), .D(CURQTDPTR1422_24), .Q(UP_DW3[24]), 
        .QN(n2568) );
    zdffb CURQTDPTR_reg_23 ( .CK(PCICLK), .D(CURQTDPTR1422_23), .Q(UP_DW3[23]), 
        .QN(n2572) );
    zdffb CURQTDPTR_reg_22 ( .CK(PCICLK), .D(CURQTDPTR1422_22), .Q(UP_DW3[22]), 
        .QN(n2576) );
    zdffb CURQTDPTR_reg_21 ( .CK(PCICLK), .D(CURQTDPTR1422_21), .Q(UP_DW3[21]), 
        .QN(n2580) );
    zdffb CURQTDPTR_reg_20 ( .CK(PCICLK), .D(CURQTDPTR1422_20), .Q(UP_DW3[20]), 
        .QN(n2584) );
    zdffb CURQTDPTR_reg_19 ( .CK(PCICLK), .D(CURQTDPTR1422_19), .Q(UP_DW3[19]), 
        .QN(n2588) );
    zdffb CURQTDPTR_reg_18 ( .CK(PCICLK), .D(CURQTDPTR1422_18), .Q(UP_DW3[18]), 
        .QN(n2592) );
    zdffb CURQTDPTR_reg_17 ( .CK(PCICLK), .D(CURQTDPTR1422_17), .Q(UP_DW3[17]), 
        .QN(n2596) );
    zdffb CURQTDPTR_reg_16 ( .CK(PCICLK), .D(CURQTDPTR1422_16), .Q(UP_DW3[16]), 
        .QN(n2600) );
    zdffb CURQTDPTR_reg_15 ( .CK(PCICLK), .D(CURQTDPTR1422_15), .Q(UP_DW3[15]), 
        .QN(n2604) );
    zdffb CURQTDPTR_reg_14 ( .CK(PCICLK), .D(CURQTDPTR1422_14), .Q(UP_DW3[14]), 
        .QN(n2608) );
    zdffb CURQTDPTR_reg_13 ( .CK(PCICLK), .D(CURQTDPTR1422_13), .Q(UP_DW3[13]), 
        .QN(n2612) );
    zdffb CURQTDPTR_reg_12 ( .CK(PCICLK), .D(CURQTDPTR1422_12), .Q(UP_DW3[12]), 
        .QN(n2616) );
    zdffb CURQTDPTR_reg_11 ( .CK(PCICLK), .D(CURQTDPTR1422_11), .Q(UP_DW3[11]), 
        .QN(n2620) );
    zdffb CURQTDPTR_reg_10 ( .CK(PCICLK), .D(CURQTDPTR1422_10), .Q(UP_DW3[10]), 
        .QN(n2624) );
    zdffb CURQTDPTR_reg_9 ( .CK(PCICLK), .D(CURQTDPTR1422_9), .Q(UP_DW3[9]), 
        .QN(n2628) );
    zdffb CURQTDPTR_reg_8 ( .CK(PCICLK), .D(CURQTDPTR1422_8), .Q(UP_DW3[8]), 
        .QN(n2632) );
    zdffb CURQTDPTR_reg_7 ( .CK(PCICLK), .D(CURQTDPTR1422_7), .Q(UP_DW3[7]), 
        .QN(n2636) );
    zdffb CURQTDPTR_reg_6 ( .CK(PCICLK), .D(CURQTDPTR1422_6), .Q(UP_DW3[6]), 
        .QN(n2640) );
    zdffb CURQTDPTR_reg_5 ( .CK(PCICLK), .D(CURQTDPTR1422_5), .Q(UP_DW3[5]), 
        .QN(n2644) );
    zdffqrb QHSM_reg_9 ( .CK(PCICLK), .D(n2286), .R(TRST_), .Q(QHSM[9]) );
    zivb U1445 ( .A(QHSM[9]), .Y(n2970) );
    zdffqrb QHSM_reg_13 ( .CK(PCICLK), .D(QHSMNXT_13), .R(TRST_), .Q(QHSM[13])
         );
    zivb U1446 ( .A(QHSM[13]), .Y(n3059) );
    zdffqrb PARSEQHEND_reg ( .CK(PCICLK), .D(PARSEQHEND_PRE), .R(TRST_), .Q(
        PARSEQHEND) );
    zdffqrb QEOT_reg ( .CK(PCICLK), .D(QEOT1815), .R(TRST_), .Q(QEOT) );
    zdffqrb_ UP_CACHE1_reg ( .CK(PCICLK), .D(QHSM[2]), .R(TRST_), .Q(UP_LDW3)
         );
    zdffqrb SPLITXSTATE_reg ( .CK(PCICLK), .D(SPLITXSTATE1256), .R(TRST_), .Q(
        TRAN_CMD[14]) );
    zivb U1447 ( .A(TRAN_CMD[14]), .Y(n2910) );
    zdffqrb QHSM_reg_7 ( .CK(PCICLK), .D(QHSMNXT_7), .R(TRST_), .Q(QHSM[7]) );
    zivb U1448 ( .A(QHSM[7]), .Y(n3048) );
    zdffb ACTIVE_reg ( .CK(PCICLK), .D(ACTIVE_NXT), .Q(ACTIVE), .QN(n2959) );
    zdffqrb QHSM_reg_6 ( .CK(PCICLK), .D(n2287), .R(TRST_), .Q(QHSM[6]) );
    zivb U1449 ( .A(QHSM[6]), .Y(n2974) );
    zdffqrb QHSM_reg_8 ( .CK(PCICLK), .D(n2285), .R(TRST_), .Q(QHSM[8]) );
    zivb U1450 ( .A(QHSM[8]), .Y(n3047) );
    zdffrb PING_ERR_reg ( .CK(PCICLK), .D(PING_ERR783), .R(TRST_), .Q(UP_DW6
        [0]), .QN(n2939) );
    zdffqrb IMMEDRETRY_reg ( .CK(PCICLK), .D(IMMEDRETRY1293), .R(TRST_), .Q(
        IMMEDRETRY) );
    zivb U1451 ( .A(IMMEDRETRY), .Y(n3052) );
    zdffqrb QHSM_reg_1 ( .CK(PCICLK), .D(QHSMNXT_1), .R(TRST_), .Q(QHSM[1]) );
    zivb U1452 ( .A(QHSM[1]), .Y(n2942) );
    zdffqrb ASYNC_EMPTY_reg ( .CK(PCICLK), .D(ASYNC_EMPTY1852), .R(TRST_), .Q(
        ASYNC_EMPTY) );
    zdffqrb_ QRXERR_CUR_reg ( .CK(PCICLK), .D(QRXERR_CUR1331), .R(TRST_), .Q(
        QRXERR) );
    zdffb XACTERR_reg ( .CK(PCICLK), .D(XACTERR1233), .QN(n2901) );
    zdffqrb_ UP_CACHE2_reg ( .CK(PCICLK), .D(QHSM[11]), .R(TRST_), .Q(UP_LDW7)
         );
    zdffqrb QHSM_reg_10 ( .CK(PCICLK), .D(QHSMNXT_10), .R(TRST_), .Q(QHSM[10])
         );
    zivb U1453 ( .A(QHSM[10]), .Y(n2977) );
    zdffqrb CACHE_INVALID_reg ( .CK(PCICLK), .D(CACHE_INVALID1602), .R(TRST_), 
        .Q(CACHE_INVALID) );
    zdffqrb CACHE_MODIFY_reg ( .CK(PCICLK), .D(CACHE_MODIFY497), .R(TRST_), 
        .Q(CACHE_MODIFY) );
    zdffqrb QHIOCINT_T_reg ( .CK(EHCIFLOW_PCLK), .D(QHIOCINT_T1889), .R(TRST_), 
        .Q(QHIOCINT_T) );
    zivb U1454 ( .A(QHIOCINT_T), .Y(n2647) );
    zdffqrb QHSM_reg_4 ( .CK(PCICLK), .D(QHSMNXT_4), .R(TRST_), .Q(QHSM[4]) );
    zivb U1455 ( .A(QHSM[4]), .Y(n3053) );
    zdffqrb QHSM_reg_5 ( .CK(PCICLK), .D(QHSMNXT_5), .R(TRST_), .Q(QHSM[5]) );
    zivb U1456 ( .A(QHSM[5]), .Y(n3055) );
    zdffqrb QCMDSTART_EOT_reg ( .CK(PCICLK), .D(QCMDSTART_EOT1778), .R(TRST_), 
        .Q(QCMDSTART_EOT) );
    zivb U1457 ( .A(QCMDSTART_EOT), .Y(n2509) );
    zdffqrb QHERRINT_reg ( .CK(EHCIFLOW_PCLK), .D(QHERRINT2000), .R(TRST_), 
        .Q(QHERRINT) );
    zdffqrb QHIOCINT_reg ( .CK(EHCIFLOW_PCLK), .D(QHIOCINT1926), .R(TRST_), 
        .Q(QHIOCINT) );
    zdffqrb QHSM_reg_11 ( .CK(PCICLK), .D(PHASENXT_resultwb), .R(TRST_), .Q(
        QHSM[11]) );
    zivb U1458 ( .A(QHSM[11]), .Y(n3051) );
    zdffqrb QHERRINT_T_reg ( .CK(EHCIFLOW_PCLK), .D(QHERRINT_T1963), .R(TRST_), 
        .Q(QHERRINT_T) );
    zivb U1459 ( .A(QHERRINT_T), .Y(n2531) );
    zdffqb QTDHALT_reg ( .CK(PCICLK), .D(n2314), .Q(QTDHALT) );
    zivb U1460 ( .A(QTDHALT), .Y(n3095) );
    zdffqb DT_reg ( .CK(PCICLK), .D(DT881), .Q(UP_DW6[31]) );
    zivb U1461 ( .A(UP_DW6[31]), .Y(n2516) );
    zivc U1462 ( .A(n3187), .Y(QHDWNUM[0]) );
    zdffrb TOTALBYTES_reg_12 ( .CK(PCICLK), .D(TOTALBYTES640_12), .R(TRST_), 
        .Q(TOTALBYTES_12), .QN(n2428) );
    zdffrb TOTALBYTES_reg_11 ( .CK(PCICLK), .D(TOTALBYTES640_11), .R(TRST_), 
        .Q(TOTALBYTES_11), .QN(n2429) );
    zdffb CERR_reg_1 ( .CK(PCICLK), .D(CERR1176_1), .Q(CERR_1), .QN(n2490) );
    znr2b U1463 ( .A(n2325), .B(n2912), .Y(n2285) );
    znr3b U1464 ( .A(GEN_PERR), .B(n2913), .C(n2975), .Y(n2286) );
    znr2b U1465 ( .A(n2325), .B(n2915), .Y(n2287) );
    znr2b U1466 ( .A(RECLAMATION), .B(n2967), .Y(n2288) );
    znr2b U1467 ( .A(n2534), .B(n2652), .Y(n2289) );
    znr3d U1468 ( .A(QH_PARSE_GO), .B(n3082), .C(n2652), .Y(n2290) );
    znr3d U1469 ( .A(QH_PARSE_GO), .B(n3086), .C(n2652), .Y(n2291) );
    znr4b U1470 ( .A(QHSM[2]), .B(n2942), .C(n2927), .D(n2966), .Y(n2292) );
    znr3b U1471 ( .A(QHSM[0]), .B(n3049), .C(n2968), .Y(n2293) );
    znr5b U1472 ( .A(QHSM[10]), .B(QHSM[2]), .C(n3051), .D(n2976), .E(QHCIREQ), 
        .Y(n2294) );
    znr3d U1473 ( .A(QHSM[13]), .B(QHDWNUM[0]), .C(n3058), .Y(n2295) );
    znr3d U1474 ( .A(n2358), .B(n3059), .C(n3058), .Y(n2296) );
    znr5b U1475 ( .A(GEN_PERR), .B(DW6[6]), .C(n2288), .D(n2969), .E(n2534), 
        .Y(n2297) );
    znr3b U1476 ( .A(n3054), .B(n2514), .C(GEN_PERR), .Y(n2298) );
    znr2b U1477 ( .A(CERR_1), .B(n3046), .Y(n2299) );
    znr2b U1478 ( .A(n2662), .B(n3092), .Y(n2300) );
    znr2b U1479 ( .A(n3091), .B(n2662), .Y(n2301) );
    znr6b U1480 ( .A(RXPIDERR), .B(TOGMATCH), .C(n2979), .D(RXSTALL), .E(RXACK
        ), .F(TRAN_CMD[6]), .Y(n2302) );
    zmux21hb U1481 ( .A(TOTALBYTES_10), .B(DW1[26]), .S(LENGTMAX), .Y(MAXLEN
        [10]) );
    zmux21hb U1482 ( .A(TOTALBYTES_9), .B(DW1[25]), .S(LENGTMAX), .Y(MAXLEN[9]
        ) );
    zmux21hb U1483 ( .A(TOTALBYTES_8), .B(DW1[24]), .S(LENGTMAX), .Y(MAXLEN[8]
        ) );
    zmux21hb U1484 ( .A(TOTALBYTES_7), .B(DW1[23]), .S(LENGTMAX), .Y(MAXLEN[7]
        ) );
    zmux21hb U1485 ( .A(TOTALBYTES_6), .B(DW1[22]), .S(LENGTMAX), .Y(MAXLEN[6]
        ) );
    zmux21hb U1486 ( .A(TOTALBYTES_5), .B(DW1[21]), .S(LENGTMAX), .Y(MAXLEN[5]
        ) );
    zmux21hb U1487 ( .A(TOTALBYTES_4), .B(DW1[20]), .S(LENGTMAX), .Y(MAXLEN[4]
        ) );
    zmux21hb U1488 ( .A(TOTALBYTES_3), .B(DW1[19]), .S(LENGTMAX), .Y(MAXLEN[3]
        ) );
    zmux21hb U1489 ( .A(TOTALBYTES_2), .B(DW1[18]), .S(LENGTMAX), .Y(MAXLEN[2]
        ) );
    zmux21hb U1490 ( .A(TOTALBYTES_1), .B(DW1[17]), .S(LENGTMAX), .Y(MAXLEN[1]
        ) );
    zmux21hb U1491 ( .A(TOTALBYTES_0), .B(DW1[16]), .S(LENGTMAX), .Y(MAXLEN[0]
        ) );
    zmux21hb U1492 ( .A(DW6[6]), .B(n3096), .S(n2320), .Y(n2314) );
    zdffqb CERR_reg_0 ( .CK(PCICLK), .D(CERR1176_0), .Q(CERR_0) );
    zivb U1493 ( .A(CERR_0), .Y(n3045) );
    zmux21lb U1494 ( .A(MAXLEN[2]), .B(ACTLEN[2]), .S(n2069), .Y(n2315) );
    zmux21lb U1495 ( .A(MAXLEN[0]), .B(ACTLEN[0]), .S(n2069), .Y(n2316) );
    zmux21lb U1496 ( .A(MAXLEN[1]), .B(ACTLEN[1]), .S(n2069), .Y(n2317) );
    zivb U1497 ( .A(CPAGE_0), .Y(n3016) );
    zdffqrb TOTALBYTES_reg_2 ( .CK(PCICLK), .D(TOTALBYTES640_2), .R(TRST_), 
        .Q(TOTALBYTES_2) );
    zivb U1498 ( .A(TOTALBYTES_2), .Y(n3006) );
    zdffqrb TOTALBYTES_reg_4 ( .CK(PCICLK), .D(TOTALBYTES640_4), .R(TRST_), 
        .Q(TOTALBYTES_4) );
    zivb U1499 ( .A(TOTALBYTES_4), .Y(n3002) );
    zdffqrb TOTALBYTES_reg_3 ( .CK(PCICLK), .D(TOTALBYTES640_3), .R(TRST_), 
        .Q(TOTALBYTES_3) );
    zivb U1500 ( .A(TOTALBYTES_3), .Y(n3004) );
    zdffqrb TOTALBYTES_reg_6 ( .CK(PCICLK), .D(TOTALBYTES640_6), .R(TRST_), 
        .Q(TOTALBYTES_6) );
    zivb U1501 ( .A(TOTALBYTES_6), .Y(n2998) );
    zdffqrb TOTALBYTES_reg_5 ( .CK(PCICLK), .D(TOTALBYTES640_5), .R(TRST_), 
        .Q(TOTALBYTES_5) );
    zivb U1502 ( .A(TOTALBYTES_5), .Y(n3000) );
    zdffqrb TOTALBYTES_reg_8 ( .CK(PCICLK), .D(TOTALBYTES640_8), .R(TRST_), 
        .Q(TOTALBYTES_8) );
    zivb U1503 ( .A(TOTALBYTES_8), .Y(n2994) );
    zdffqrb TOTALBYTES_reg_7 ( .CK(PCICLK), .D(TOTALBYTES640_7), .R(TRST_), 
        .Q(TOTALBYTES_7) );
    zivb U1504 ( .A(TOTALBYTES_7), .Y(n2996) );
    zdffqrb TOTALBYTES_reg_9 ( .CK(PCICLK), .D(TOTALBYTES640_9), .R(TRST_), 
        .Q(TOTALBYTES_9) );
    zivb U1505 ( .A(TOTALBYTES_9), .Y(n2992) );
    zor2b U1506 ( .A(n2461), .B(n2459), .Y(n2318) );
    znr2b U1507 ( .A(sub_383_carry_14), .B(TOTALBYTES_14), .Y(n2319) );
    ziv11b U1508 ( .A(PHASENXT_exechk), .Y(n2320), .Z(n2321) );
    zivf U1509 ( .A(n2322), .Y(QHDWNUM[3]) );
    zivc U1510 ( .A(QHDWNUM[0]), .Y(QHSM[12]) );
    zivb U1511 ( .A(n3187), .Y(n2322) );
    zivb U1512 ( .A(n2322), .Y(n2358) );
    zivb U1513 ( .A(QHDWNUM[0]), .Y(QHCIADR[2]) );
    zoai2x4b U1514 ( .A(n2591), .B(n3159), .C(n3160), .D(n2592), .E(n2593), 
        .F(n3162), .G(n2594), .H(n3164), .Y(CURQTDPTR1422_18) );
    zoai2x4b U1515 ( .A(n2635), .B(n3159), .C(n2537), .D(n2636), .E(n2637), 
        .F(n3161), .G(n2638), .H(n3164), .Y(CURQTDPTR1422_7) );
    zoai2x4b U1516 ( .A(n2579), .B(n3159), .C(n3160), .D(n2580), .E(n2581), 
        .F(n3162), .G(n2582), .H(n3164), .Y(CURQTDPTR1422_21) );
    zoai2x4b U1517 ( .A(n2615), .B(n3159), .C(n3160), .D(n2616), .E(n2617), 
        .F(n3162), .G(n2618), .H(n3164), .Y(CURQTDPTR1422_12) );
    zoai2x4b U1518 ( .A(n2563), .B(n3159), .C(n2537), .D(n2564), .E(n2565), 
        .F(n3161), .G(n2566), .H(n3163), .Y(CURQTDPTR1422_25) );
    zoai2x4b U1519 ( .A(n2627), .B(n3159), .C(n2537), .D(n2628), .E(n2629), 
        .F(n3162), .G(n2630), .H(n3163), .Y(CURQTDPTR1422_9) );
    zor3d U1520 ( .A(n2534), .B(n2650), .C(n3090), .Y(n3159) );
    zoai2x4b U1521 ( .A(n2595), .B(n2536), .C(n2537), .D(n2596), .E(n2597), 
        .F(n2540), .G(n2598), .H(n2542), .Y(CURQTDPTR1422_17) );
    zoai2x4b U1522 ( .A(n2547), .B(n2536), .C(n2537), .D(n2548), .E(n2549), 
        .F(n2540), .G(n2550), .H(n2542), .Y(CURQTDPTR1422_29) );
    zoai2x4b U1523 ( .A(n2607), .B(n2536), .C(n3160), .D(n2608), .E(n2609), 
        .F(n2540), .G(n2610), .H(n2542), .Y(CURQTDPTR1422_14) );
    zoai2x4b U1524 ( .A(n2571), .B(n2536), .C(n3160), .D(n2572), .E(n2573), 
        .F(n2540), .G(n2574), .H(n2542), .Y(CURQTDPTR1422_23) );
    zoai2x4b U1525 ( .A(n2619), .B(n2536), .C(n2537), .D(n2620), .E(n2621), 
        .F(n2540), .G(n2622), .H(n2542), .Y(CURQTDPTR1422_11) );
    zoai2x4b U1526 ( .A(n2559), .B(n2536), .C(n3160), .D(n2560), .E(n2561), 
        .F(n2540), .G(n2562), .H(n2542), .Y(CURQTDPTR1422_26) );
    zor3d U1527 ( .A(n2534), .B(n2650), .C(n3090), .Y(n2536) );
    zoai2x4b U1528 ( .A(n2587), .B(n3158), .C(n2537), .D(n2588), .E(n2589), 
        .F(n3161), .G(n2590), .H(n3163), .Y(CURQTDPTR1422_19) );
    zoai2x4b U1529 ( .A(n2639), .B(n3158), .C(n3160), .D(n2640), .E(n2641), 
        .F(n3162), .G(n2642), .H(n3163), .Y(CURQTDPTR1422_6) );
    zoai2x4b U1530 ( .A(n2575), .B(n3158), .C(n2537), .D(n2576), .E(n2577), 
        .F(n3161), .G(n2578), .H(n3163), .Y(CURQTDPTR1422_22) );
    zoai2x4b U1531 ( .A(n2611), .B(n3158), .C(n2537), .D(n2612), .E(n2613), 
        .F(n3161), .G(n2614), .H(n3163), .Y(CURQTDPTR1422_13) );
    zoai2x4b U1532 ( .A(n2567), .B(n3158), .C(n2537), .D(n2568), .E(n2569), 
        .F(n3162), .G(n2570), .H(n3164), .Y(CURQTDPTR1422_24) );
    zoai2x4b U1533 ( .A(n2623), .B(n3158), .C(n3160), .D(n2624), .E(n2625), 
        .F(n3161), .G(n2626), .H(n3164), .Y(CURQTDPTR1422_10) );
    zor3d U1534 ( .A(n2534), .B(n2650), .C(n3090), .Y(n3158) );
    zivb U1535 ( .A(n3074), .Y(n2323) );
    zivd U1536 ( .A(DWCNT[1]), .Y(n3074) );
    zivb U1537 ( .A(n3070), .Y(n2324) );
    zivd U1538 ( .A(DWCNT[2]), .Y(n3070) );
    zivb U1539 ( .A(n2498), .Y(n2325) );
    zor2b U1540 ( .A(GEN_PERR), .B(n3097), .Y(n2518) );
    zor2b U1541 ( .A(GEN_PERR), .B(n2890), .Y(n2931) );
    zivc U1542 ( .A(GEN_PERR), .Y(n2498) );
    zoa21b U1543 ( .A(n2321), .B(QHSM[3]), .C(n2947), .Y(n2946) );
    zdffqrb QHSM_reg_3 ( .CK(PCICLK), .D(n2321), .R(TRST_), .Q(QHSM[3]) );
    zor2b U1544 ( .A(PHASENXT_exechk), .B(n3030), .Y(n3029) );
    zor3d U1545 ( .A(CPAGE_1), .B(CPAGE_0), .C(n2328), .Y(n2326) );
    zor3d U1546 ( .A(CPAGE_1), .B(CPAGE_0), .C(n2328), .Y(n2804) );
    zbfd U1547 ( .A(CPAGE_2), .Y(n2327) );
    zbfd U1548 ( .A(CPAGE_2), .Y(n2328) );
    zivb U1549 ( .A(n2328), .Y(n3012) );
    zdffqb CPAGE_reg_2 ( .CK(PCICLK), .D(CPAGE1098_2), .Q(CPAGE_2) );
    zbfb U1550 ( .A(DW1[12]), .Y(TRAN_CMD[13]) );
    zbfb U1551 ( .A(DW2[23]), .Y(TRAN_CMD[15]) );
    zbfb U1552 ( .A(DW2[24]), .Y(TRAN_CMD[16]) );
    zbfb U1553 ( .A(DW2[25]), .Y(TRAN_CMD[17]) );
    zbfb U1554 ( .A(DW2[26]), .Y(TRAN_CMD[18]) );
    zbfb U1555 ( .A(DW2[27]), .Y(TRAN_CMD[19]) );
    zbfb U1556 ( .A(DW2[28]), .Y(TRAN_CMD[20]) );
    zbfb U1557 ( .A(DW2[29]), .Y(TRAN_CMD[21]) );
    zbfb U1558 ( .A(DW2[16]), .Y(TRAN_CMD[22]) );
    zbfb U1559 ( .A(DW2[17]), .Y(TRAN_CMD[23]) );
    zbfb U1560 ( .A(DW2[18]), .Y(TRAN_CMD[24]) );
    zbfb U1561 ( .A(DW2[19]), .Y(TRAN_CMD[25]) );
    zbfb U1562 ( .A(DW2[20]), .Y(TRAN_CMD[26]) );
    zbfb U1563 ( .A(DW2[21]), .Y(TRAN_CMD[27]) );
    zbfb U1564 ( .A(DW2[22]), .Y(TRAN_CMD[28]) );
    zbfb U1565 ( .A(DW1[8]), .Y(TRAN_CMD[29]) );
    zbfb U1566 ( .A(DW1[9]), .Y(TRAN_CMD[30]) );
    zbfb U1567 ( .A(DW1[10]), .Y(TRAN_CMD[31]) );
    zbfb U1568 ( .A(DW1[11]), .Y(TRAN_CMD[32]) );
    zbfb U1569 ( .A(DW1[0]), .Y(TRAN_CMD[33]) );
    zbfb U1570 ( .A(DW1[1]), .Y(TRAN_CMD[34]) );
    zbfb U1571 ( .A(DW1[2]), .Y(TRAN_CMD[35]) );
    zbfb U1572 ( .A(DW1[3]), .Y(TRAN_CMD[36]) );
    zbfb U1573 ( .A(DW1[4]), .Y(TRAN_CMD[37]) );
    zbfb U1574 ( .A(DW1[5]), .Y(TRAN_CMD[38]) );
    zbfb U1575 ( .A(DW1[6]), .Y(TRAN_CMD[39]) );
    zbfb U1576 ( .A(QHCIMWR), .Y(QHCIADR[3]) );
    zor2b U1577 ( .A(n3187), .B(QHSM[13]), .Y(QHCIMWR) );
    zbfb U1578 ( .A(QHDWNUM[2]), .Y(QHDWNUM[1]) );
    zivb U1579 ( .A(QHCIMWR), .Y(QHDWNUM[2]) );
    zdffqrb QHSM_reg_12 ( .CK(PCICLK), .D(QHSMNXT_12), .R(TRST_), .Q(n3187) );
    zbfb U1580 ( .A(UP_LDW6), .Y(UP_LDW5) );
    zor2b U1581 ( .A(UP_LDW3), .B(UP_LDW7), .Y(UP_LDW6) );
    zbfb U1582 ( .A(UP_DW7[0]), .Y(TRAN_CMD[72]) );
    zdffqb OVERWBOFFSET_reg_0 ( .CK(PCICLK), .D(OVERWBOFFSET1715_0), .Q(UP_DW7
        [0]) );
    zbfb U1583 ( .A(UP_DW7[1]), .Y(TRAN_CMD[73]) );
    zdffqb OVERWBOFFSET_reg_1 ( .CK(PCICLK), .D(OVERWBOFFSET1715_1), .Q(UP_DW7
        [1]) );
    zbfb U1584 ( .A(UP_DW7[2]), .Y(TRAN_CMD[74]) );
    zdffqb OVERWBOFFSET_reg_2 ( .CK(PCICLK), .D(OVERWBOFFSET1715_2), .Q(UP_DW7
        [2]) );
    zbfb U1585 ( .A(UP_DW7[3]), .Y(TRAN_CMD[75]) );
    zdffqb OVERWBOFFSET_reg_3 ( .CK(PCICLK), .D(OVERWBOFFSET1715_3), .Q(UP_DW7
        [3]) );
    zbfb U1586 ( .A(UP_DW7[4]), .Y(TRAN_CMD[76]) );
    zdffqb OVERWBOFFSET_reg_4 ( .CK(PCICLK), .D(OVERWBOFFSET1715_4), .Q(UP_DW7
        [4]) );
    zbfb U1587 ( .A(UP_DW7[5]), .Y(TRAN_CMD[77]) );
    zdffqb OVERWBOFFSET_reg_5 ( .CK(PCICLK), .D(OVERWBOFFSET1715_5), .Q(UP_DW7
        [5]) );
    zbfb U1588 ( .A(UP_DW7[6]), .Y(TRAN_CMD[78]) );
    zdffqb OVERWBOFFSET_reg_6 ( .CK(PCICLK), .D(OVERWBOFFSET1715_6), .Q(UP_DW7
        [6]) );
    zbfb U1589 ( .A(UP_DW7[7]), .Y(TRAN_CMD[79]) );
    zdffqb OVERWBOFFSET_reg_7 ( .CK(PCICLK), .D(OVERWBOFFSET1715_7), .Q(UP_DW7
        [7]) );
    zbfb U1590 ( .A(UP_DW7[8]), .Y(TRAN_CMD[80]) );
    zdffqb OVERWBOFFSET_reg_8 ( .CK(PCICLK), .D(OVERWBOFFSET1715_8), .Q(UP_DW7
        [8]) );
    zbfb U1591 ( .A(UP_DW7[9]), .Y(TRAN_CMD[81]) );
    zdffqb OVERWBOFFSET_reg_9 ( .CK(PCICLK), .D(OVERWBOFFSET1715_9), .Q(UP_DW7
        [9]) );
    zbfb U1592 ( .A(UP_DW7[10]), .Y(TRAN_CMD[82]) );
    zdffqb OVERWBOFFSET_reg_10 ( .CK(PCICLK), .D(OVERWBOFFSET1715_10), .Q(
        UP_DW7[10]) );
    zbfb U1593 ( .A(UP_DW7[11]), .Y(TRAN_CMD[83]) );
    zdffqb OVERWBOFFSET_reg_11 ( .CK(PCICLK), .D(OVERWBOFFSET1715_11), .Q(
        UP_DW7[11]) );
    zbfb U1594 ( .A(DW7[12]), .Y(UP_DW7[12]) );
    zbfb U1595 ( .A(DW7[13]), .Y(UP_DW7[13]) );
    zbfb U1596 ( .A(DW7[14]), .Y(UP_DW7[14]) );
    zbfb U1597 ( .A(DW7[15]), .Y(UP_DW7[15]) );
    zbfb U1598 ( .A(DW7[16]), .Y(UP_DW7[16]) );
    zbfb U1599 ( .A(DW7[17]), .Y(UP_DW7[17]) );
    zbfb U1600 ( .A(DW7[18]), .Y(UP_DW7[18]) );
    zbfb U1601 ( .A(DW7[19]), .Y(UP_DW7[19]) );
    zbfb U1602 ( .A(DW7[20]), .Y(UP_DW7[20]) );
    zbfb U1603 ( .A(DW7[21]), .Y(UP_DW7[21]) );
    zbfb U1604 ( .A(DW7[22]), .Y(UP_DW7[22]) );
    zbfb U1605 ( .A(DW7[23]), .Y(UP_DW7[23]) );
    zbfb U1606 ( .A(DW7[24]), .Y(UP_DW7[24]) );
    zbfb U1607 ( .A(DW7[25]), .Y(UP_DW7[25]) );
    zbfb U1608 ( .A(DW7[26]), .Y(UP_DW7[26]) );
    zbfb U1609 ( .A(DW7[27]), .Y(UP_DW7[27]) );
    zbfb U1610 ( .A(DW7[28]), .Y(UP_DW7[28]) );
    zbfb U1611 ( .A(DW7[29]), .Y(UP_DW7[29]) );
    zbfb U1612 ( .A(DW7[30]), .Y(UP_DW7[30]) );
    zbfb U1613 ( .A(DW7[31]), .Y(UP_DW7[31]) );
    zbfb U1614 ( .A(DW6[9]), .Y(UP_DW6[9]) );
    zbfb U1615 ( .A(DW6[15]), .Y(UP_DW6[15]) );
    zbfb U1616 ( .A(DW5[0]), .Y(UP_DW5[0]) );
    zbfb U1617 ( .A(DW5[5]), .Y(UP_DW5[5]) );
    zbfb U1618 ( .A(DW5[6]), .Y(UP_DW5[6]) );
    zbfb U1619 ( .A(DW5[7]), .Y(UP_DW5[7]) );
    zbfb U1620 ( .A(DW5[8]), .Y(UP_DW5[8]) );
    zbfb U1621 ( .A(DW5[9]), .Y(UP_DW5[9]) );
    zbfb U1622 ( .A(DW5[10]), .Y(UP_DW5[10]) );
    zbfb U1623 ( .A(DW5[11]), .Y(UP_DW5[11]) );
    zbfb U1624 ( .A(DW5[12]), .Y(UP_DW5[12]) );
    zbfb U1625 ( .A(DW5[13]), .Y(UP_DW5[13]) );
    zbfb U1626 ( .A(DW5[14]), .Y(UP_DW5[14]) );
    zbfb U1627 ( .A(DW5[15]), .Y(UP_DW5[15]) );
    zbfb U1628 ( .A(DW5[16]), .Y(UP_DW5[16]) );
    zbfb U1629 ( .A(DW5[17]), .Y(UP_DW5[17]) );
    zbfb U1630 ( .A(DW5[18]), .Y(UP_DW5[18]) );
    zbfb U1631 ( .A(DW5[19]), .Y(UP_DW5[19]) );
    zbfb U1632 ( .A(DW5[20]), .Y(UP_DW5[20]) );
    zbfb U1633 ( .A(DW5[21]), .Y(UP_DW5[21]) );
    zbfb U1634 ( .A(DW5[22]), .Y(UP_DW5[22]) );
    zbfb U1635 ( .A(DW5[23]), .Y(UP_DW5[23]) );
    zbfb U1636 ( .A(DW5[24]), .Y(UP_DW5[24]) );
    zbfb U1637 ( .A(DW5[25]), .Y(UP_DW5[25]) );
    zbfb U1638 ( .A(DW5[26]), .Y(UP_DW5[26]) );
    zbfb U1639 ( .A(DW5[27]), .Y(UP_DW5[27]) );
    zbfb U1640 ( .A(DW5[28]), .Y(UP_DW5[28]) );
    zbfb U1641 ( .A(DW5[29]), .Y(UP_DW5[29]) );
    zbfb U1642 ( .A(DW5[30]), .Y(UP_DW5[30]) );
    zbfb U1643 ( .A(DW5[31]), .Y(UP_DW5[31]) );
    zbfb U1644 ( .A(QHSM[0]), .Y(QHIDLE) );
    zdffqsb QHSM_reg_0 ( .CK(PCICLK), .D(PHASENXT_idle), .S(TRST_), .Q(QHSM[0]
        ) );
    zan2b U1645 ( .A(UP_DW7[11]), .B(r285_carry_11), .Y(OVERWBOFFSET_P1671_12)
         );
    zxo2b U1646 ( .A(UP_DW7[11]), .B(r285_carry_11), .Y(OVERWBOFFSET_P1671_11)
         );
    zan2b U1647 ( .A(_cell_705_U89_Z_0), .B(UP_DW7[0]), .Y(r285_carry_1) );
    zxo2b U1648 ( .A(_cell_705_U89_Z_0), .B(UP_DW7[0]), .Y(
        OVERWBOFFSET_P1671_0) );
    zxn2b U1649 ( .A(sub_383_carry_14), .B(TOTALBYTES_14), .Y(
        VIR_TOTALBYTES_14) );
    zor2b U1650 ( .A(sub_383_carry_13), .B(TOTALBYTES_13), .Y(sub_383_carry_14
        ) );
    zxn2b U1651 ( .A(sub_383_carry_13), .B(TOTALBYTES_13), .Y(
        VIR_TOTALBYTES_13) );
    zor2b U1652 ( .A(sub_383_carry_12), .B(TOTALBYTES_12), .Y(sub_383_carry_13
        ) );
    zxn2b U1653 ( .A(sub_383_carry_12), .B(TOTALBYTES_12), .Y(
        VIR_TOTALBYTES_12) );
    zor2b U1654 ( .A(sub_383_carry_11), .B(TOTALBYTES_11), .Y(sub_383_carry_12
        ) );
    zxn2b U1655 ( .A(sub_383_carry_11), .B(TOTALBYTES_11), .Y(
        VIR_TOTALBYTES_11) );
    zor2b U1656 ( .A(TOTALBYTES_0), .B(n2316), .Y(sub_383_carry_1) );
    zxn2b U1657 ( .A(TOTALBYTES_0), .B(n2316), .Y(VIR_TOTALBYTES_0) );
    zymx24hb U1658 ( .A1(MAXLEN[6]), .A2(MAXLEN[5]), .A3(MAXLEN[4]), .A4(
        MAXLEN[3]), .B1(ACTLEN[6]), .B2(ACTLEN[5]), .B3(ACTLEN[4]), .B4(ACTLEN
        [3]), .S(n2069), .Y1(MINUEND_6), .Y2(MINUEND_5), .Y3(MINUEND_4), .Y4(
        MINUEND_3) );
    zymx24hb U1659 ( .A1(MAXLEN[10]), .A2(MAXLEN[9]), .A3(MAXLEN[8]), .A4(
        MAXLEN[7]), .B1(ACTLEN[10]), .B2(ACTLEN[9]), .B3(ACTLEN[8]), .B4(
        ACTLEN[7]), .S(n2069), .Y1(MINUEND_10), .Y2(MINUEND_9), .Y3(MINUEND_8), 
        .Y4(MINUEND_7) );
    zdffqd CPAGE_reg_1 ( .CK(PCICLK), .D(CPAGE1098_1), .Q(CPAGE_1) );
    zdffqd CPAGE_reg_0 ( .CK(PCICLK), .D(CPAGE1098_0), .Q(CPAGE_0) );
    zdffqrd QHSM_reg_2 ( .CK(PCICLK), .D(QHSMNXT_2), .R(TRST_), .Q(QHSM[2]) );
    znd2d U1660 ( .A(n2482), .B(n2318), .Y(LENGTMAX) );
    zfa1b sub_383_U2_6 ( .A(TOTALBYTES_6), .B(sub_383_B_not_6), .CI(
        sub_383_carry_6), .CO(sub_383_carry_7), .S(VIR_TOTALBYTES_6) );
    zfa1b sub_383_U2_8 ( .A(TOTALBYTES_8), .B(sub_383_B_not_8), .CI(
        sub_383_carry_8), .CO(sub_383_carry_9), .S(VIR_TOTALBYTES_8) );
    zfa1b sub_383_U2_10 ( .A(TOTALBYTES_10), .B(sub_383_B_not_10), .CI(
        sub_383_carry_10), .CO(sub_383_carry_11), .S(VIR_TOTALBYTES_10) );
    zfa1b sub_383_U2_9 ( .A(TOTALBYTES_9), .B(sub_383_B_not_9), .CI(
        sub_383_carry_9), .CO(sub_383_carry_10), .S(VIR_TOTALBYTES_9) );
    zfa1b sub_383_U2_1 ( .A(TOTALBYTES_1), .B(n2317), .CI(sub_383_carry_1), 
        .CO(sub_383_carry_2), .S(VIR_TOTALBYTES_1) );
    zfa1b sub_383_U2_7 ( .A(TOTALBYTES_7), .B(sub_383_B_not_7), .CI(
        sub_383_carry_7), .CO(sub_383_carry_8), .S(VIR_TOTALBYTES_7) );
    zfa1b sub_383_U2_5 ( .A(TOTALBYTES_5), .B(sub_383_B_not_5), .CI(
        sub_383_carry_5), .CO(sub_383_carry_6), .S(VIR_TOTALBYTES_5) );
    zfa1b sub_383_U2_3 ( .A(TOTALBYTES_3), .B(sub_383_B_not_3), .CI(
        sub_383_carry_3), .CO(sub_383_carry_4), .S(VIR_TOTALBYTES_3) );
    zfa1b sub_383_U2_2 ( .A(TOTALBYTES_2), .B(n2315), .CI(sub_383_carry_2), 
        .CO(sub_383_carry_3), .S(VIR_TOTALBYTES_2) );
    zfa1b sub_383_U2_4 ( .A(TOTALBYTES_4), .B(sub_383_B_not_4), .CI(
        sub_383_carry_4), .CO(sub_383_carry_5), .S(VIR_TOTALBYTES_4) );
    zfa1b r285_U1_5 ( .A(UP_DW7[5]), .B(_cell_705_U89_Z_5), .CI(r285_carry_5), 
        .CO(r285_carry_6), .S(OVERWBOFFSET_P1671_5) );
    zfa1b r285_U1_4 ( .A(UP_DW7[4]), .B(_cell_705_U89_Z_4), .CI(r285_carry_4), 
        .CO(r285_carry_5), .S(OVERWBOFFSET_P1671_4) );
    zfa1b r285_U1_3 ( .A(UP_DW7[3]), .B(_cell_705_U89_Z_3), .CI(r285_carry_3), 
        .CO(r285_carry_4), .S(OVERWBOFFSET_P1671_3) );
    zfa1b r285_U1_10 ( .A(UP_DW7[10]), .B(_cell_705_U89_Z_10), .CI(
        r285_carry_10), .CO(r285_carry_11), .S(OVERWBOFFSET_P1671_10) );
    zfa1b r285_U1_9 ( .A(UP_DW7[9]), .B(_cell_705_U89_Z_9), .CI(r285_carry_9), 
        .CO(r285_carry_10), .S(OVERWBOFFSET_P1671_9) );
    zfa1b r285_U1_2 ( .A(UP_DW7[2]), .B(_cell_705_U89_Z_2), .CI(r285_carry_2), 
        .CO(r285_carry_3), .S(OVERWBOFFSET_P1671_2) );
    zfa1b r285_U1_7 ( .A(UP_DW7[7]), .B(_cell_705_U89_Z_7), .CI(r285_carry_7), 
        .CO(r285_carry_8), .S(OVERWBOFFSET_P1671_7) );
    zfa1b r285_U1_8 ( .A(UP_DW7[8]), .B(_cell_705_U89_Z_8), .CI(r285_carry_8), 
        .CO(r285_carry_9), .S(OVERWBOFFSET_P1671_8) );
    zfa1b r285_U1_6 ( .A(UP_DW7[6]), .B(_cell_705_U89_Z_6), .CI(r285_carry_6), 
        .CO(r285_carry_7), .S(OVERWBOFFSET_P1671_6) );
    zfa1b r285_U1_1 ( .A(UP_DW7[1]), .B(_cell_705_U89_Z_1), .CI(r285_carry_1), 
        .CO(r285_carry_2), .S(OVERWBOFFSET_P1671_1) );
    zao211b U1661 ( .A(n2491), .B(n2492), .C(n2493), .D(n2494), .Y(
        PHASENXT_idle) );
    zind2d U1662 ( .A(DW1[12]), .B(DW1[13]), .Y(TRAN_CMD[6]) );
    zao21d U1663 ( .A(DW6[7]), .B(n2297), .C(n2495), .Y(PHASENXT_exechk) );
    zor6b U1664 ( .A(n2286), .B(n2285), .C(QHSMNXT_7), .D(QHSMNXT_4), .E(n2287
        ), .F(QHSMNXT_5), .Y(QTDEXE) );
    zoa21d U1665 ( .A(n2507), .B(n2508), .C(n2509), .Y(QCMDSTART_REQ) );
    zoa21d U1666 ( .A(QCMDSTART_EOT), .B(QCMDSTART), .C(n2514), .Y(
        QCMDSTART_EOT1778) );
    zoa21d U1667 ( .A(TRAN_CMD[7]), .B(n2516), .C(n2511), .Y(TRAN_CMD[4]) );
    zan4b U1668 ( .A(n2517), .B(n2518), .C(n2505), .D(n2519), .Y(QHPARSING) );
    zan4b U1669 ( .A(PCIEND), .B(n2292), .C(DW6[7]), .D(n2498), .Y(QHSMNXT_2)
         );
    zao222b U1671 ( .A(UP_DW7[0]), .B(n2653), .C(DW7[0]), .D(n2654), .E(
        OVERWBOFFSET_P1671_0), .F(n2655), .Y(OVERWBOFFSET1715_0) );
    zao222b U1672 ( .A(UP_DW7[1]), .B(n2653), .C(DW7[1]), .D(n2654), .E(
        OVERWBOFFSET_P1671_1), .F(n2655), .Y(OVERWBOFFSET1715_1) );
    zao222b U1673 ( .A(UP_DW7[2]), .B(n2653), .C(DW7[2]), .D(n2654), .E(
        OVERWBOFFSET_P1671_2), .F(n2655), .Y(OVERWBOFFSET1715_2) );
    zao222b U1674 ( .A(UP_DW7[3]), .B(n2653), .C(DW7[3]), .D(n2654), .E(
        OVERWBOFFSET_P1671_3), .F(n2655), .Y(OVERWBOFFSET1715_3) );
    zao222b U1675 ( .A(UP_DW7[4]), .B(n2653), .C(DW7[4]), .D(n2654), .E(
        OVERWBOFFSET_P1671_4), .F(n2655), .Y(OVERWBOFFSET1715_4) );
    zao222b U1676 ( .A(UP_DW7[5]), .B(n2653), .C(DW7[5]), .D(n2654), .E(
        OVERWBOFFSET_P1671_5), .F(n2655), .Y(OVERWBOFFSET1715_5) );
    zao222b U1677 ( .A(UP_DW7[6]), .B(n2653), .C(DW7[6]), .D(n2654), .E(
        OVERWBOFFSET_P1671_6), .F(n2655), .Y(OVERWBOFFSET1715_6) );
    zao222b U1678 ( .A(UP_DW7[7]), .B(n2653), .C(DW7[7]), .D(n2654), .E(
        OVERWBOFFSET_P1671_7), .F(n2655), .Y(OVERWBOFFSET1715_7) );
    zao222b U1679 ( .A(UP_DW7[8]), .B(n2653), .C(DW7[8]), .D(n2654), .E(
        OVERWBOFFSET_P1671_8), .F(n2655), .Y(OVERWBOFFSET1715_8) );
    zao222b U1680 ( .A(UP_DW7[9]), .B(n2653), .C(DW7[9]), .D(n2654), .E(
        OVERWBOFFSET_P1671_9), .F(n2655), .Y(OVERWBOFFSET1715_9) );
    zao222b U1681 ( .A(UP_DW7[10]), .B(n2653), .C(DW7[10]), .D(n2654), .E(
        OVERWBOFFSET_P1671_10), .F(n2655), .Y(OVERWBOFFSET1715_10) );
    zao222b U1682 ( .A(UP_DW7[11]), .B(n2653), .C(DW7[11]), .D(n2654), .E(
        OVERWBOFFSET_P1671_11), .F(n2655), .Y(OVERWBOFFSET1715_11) );
    zan4b U1683 ( .A(n2650), .B(n2497), .C(n2659), .D(n2660), .Y(
        QRXERR_CUR1331) );
    zao222b U1684 ( .A(DW6[14]), .B(n2662), .C(n2301), .D(n2328), .E(
        CPAGE1102_2), .F(n2300), .Y(CPAGE1098_2) );
    zao222b U1685 ( .A(DW6[13]), .B(n2662), .C(n2301), .D(CPAGE_1), .E(
        CPAGE1102_1), .F(n2300), .Y(CPAGE1098_1) );
    zao222b U1686 ( .A(DW6[12]), .B(n2662), .C(n2301), .D(CPAGE_0), .E(n3016), 
        .F(n2300), .Y(CPAGE1098_0) );
    zao222b U1687 ( .A(n2663), .B(TOTALBYTES_14), .C(DW6[30]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_14), .F(n2664), .Y(
        TOTALBYTES640_14) );
    zao222b U1688 ( .A(n2663), .B(TOTALBYTES_13), .C(DW6[29]), .D(n2321), .E(
        VIR_TOTALBYTES_13), .F(n2664), .Y(TOTALBYTES640_13) );
    zao222b U1689 ( .A(n2663), .B(TOTALBYTES_12), .C(DW6[28]), .D(n2321), .E(
        VIR_TOTALBYTES_12), .F(n2664), .Y(TOTALBYTES640_12) );
    zao222b U1690 ( .A(n2663), .B(TOTALBYTES_11), .C(DW6[27]), .D(n2321), .E(
        VIR_TOTALBYTES_11), .F(n2664), .Y(TOTALBYTES640_11) );
    zao222b U1691 ( .A(n2663), .B(TOTALBYTES_10), .C(DW6[26]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_10), .F(n2664), .Y(
        TOTALBYTES640_10) );
    zao222b U1692 ( .A(n2663), .B(TOTALBYTES_9), .C(DW6[25]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_9), .F(n2664), .Y(TOTALBYTES640_9)
         );
    zao222b U1693 ( .A(n2663), .B(TOTALBYTES_8), .C(DW6[24]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_8), .F(n2664), .Y(TOTALBYTES640_8)
         );
    zao222b U1694 ( .A(n2663), .B(TOTALBYTES_7), .C(DW6[23]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_7), .F(n2664), .Y(TOTALBYTES640_7)
         );
    zao222b U1695 ( .A(n2663), .B(TOTALBYTES_6), .C(DW6[22]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_6), .F(n2664), .Y(TOTALBYTES640_6)
         );
    zao222b U1696 ( .A(n2663), .B(TOTALBYTES_5), .C(DW6[21]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_5), .F(n2664), .Y(TOTALBYTES640_5)
         );
    zao222b U1697 ( .A(n2663), .B(TOTALBYTES_4), .C(DW6[20]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_4), .F(n2664), .Y(TOTALBYTES640_4)
         );
    zao222b U1698 ( .A(n2663), .B(TOTALBYTES_3), .C(DW6[19]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_3), .F(n2664), .Y(TOTALBYTES640_3)
         );
    zao222b U1699 ( .A(n2663), .B(TOTALBYTES_2), .C(DW6[18]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_2), .F(n2664), .Y(TOTALBYTES640_2)
         );
    zao222b U1700 ( .A(n2663), .B(TOTALBYTES_1), .C(DW6[17]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_1), .F(n2664), .Y(TOTALBYTES640_1)
         );
    zao222b U1701 ( .A(n2663), .B(TOTALBYTES_0), .C(DW6[16]), .D(
        PHASENXT_exechk), .E(VIR_TOTALBYTES_0), .F(n2664), .Y(TOTALBYTES640_0)
         );
    zor3b U1702 ( .A(n2665), .B(n2666), .C(n2667), .Y(QHCIADD[0]) );
    zor3b U1703 ( .A(n2668), .B(n2669), .C(n2670), .Y(QHCIADD[1]) );
    zor3b U1704 ( .A(n2671), .B(n2672), .C(n2673), .Y(QHCIADD[2]) );
    zor3b U1705 ( .A(n2674), .B(n2675), .C(n2676), .Y(QHCIADD[3]) );
    zor3b U1706 ( .A(n2677), .B(n2678), .C(n2679), .Y(QHCIADD[4]) );
    zor3b U1707 ( .A(n2680), .B(n2681), .C(n2682), .Y(QHCIADD[5]) );
    zor3b U1708 ( .A(n2683), .B(n2684), .C(n2685), .Y(QHCIADD[6]) );
    zor3b U1709 ( .A(n2686), .B(n2687), .C(n2688), .Y(QHCIADD[7]) );
    zor3b U1710 ( .A(n2689), .B(n2690), .C(n2691), .Y(QHCIADD[8]) );
    zor3b U1711 ( .A(n2692), .B(n2693), .C(n2694), .Y(QHCIADD[9]) );
    zor3b U1712 ( .A(n2695), .B(n2696), .C(n2697), .Y(QHCIADD[10]) );
    zor3b U1713 ( .A(n2698), .B(n2699), .C(n2700), .Y(QHCIADD[11]) );
    zor3b U1714 ( .A(n2701), .B(n2702), .C(n2703), .Y(QHCIADD[12]) );
    zor3b U1715 ( .A(n2704), .B(n2705), .C(n2706), .Y(QHCIADD[13]) );
    zor3b U1716 ( .A(n2707), .B(n2708), .C(n2709), .Y(QHCIADD[14]) );
    zor3b U1717 ( .A(n2710), .B(n2711), .C(n2712), .Y(QHCIADD[15]) );
    zor3b U1718 ( .A(n2713), .B(n2714), .C(n2715), .Y(QHCIADD[16]) );
    zor3b U1719 ( .A(n2716), .B(n2717), .C(n2718), .Y(QHCIADD[17]) );
    zor3b U1720 ( .A(n2719), .B(n2720), .C(n2721), .Y(QHCIADD[18]) );
    zor3b U1721 ( .A(n2722), .B(n2723), .C(n2724), .Y(QHCIADD[19]) );
    zor3b U1722 ( .A(n2725), .B(n2726), .C(n2727), .Y(QHCIADD[20]) );
    zor3b U1723 ( .A(n2728), .B(n2729), .C(n2730), .Y(QHCIADD[21]) );
    zor3b U1724 ( .A(n2731), .B(n2732), .C(n2733), .Y(QHCIADD[22]) );
    zor3b U1725 ( .A(n2734), .B(n2735), .C(n2736), .Y(QHCIADD[23]) );
    zor3b U1726 ( .A(n2737), .B(n2738), .C(n2739), .Y(QHCIADD[24]) );
    zor3b U1727 ( .A(n2740), .B(n2741), .C(n2742), .Y(QHCIADD[25]) );
    zor3b U1728 ( .A(n2743), .B(n2744), .C(n2745), .Y(QHCIADD[26]) );
    zor3b U1729 ( .A(n2746), .B(n2747), .C(n2748), .Y(QHCIADD[27]) );
    zor3b U1730 ( .A(n2749), .B(n2750), .C(n2751), .Y(QHCIADD[28]) );
    zor3b U1731 ( .A(n2752), .B(n2753), .C(n2754), .Y(QHCIADD[29]) );
    zor3b U1732 ( .A(n2755), .B(n2756), .C(n2757), .Y(QHCIADD[30]) );
    zor3b U1733 ( .A(n2758), .B(n2759), .C(n2760), .Y(QHCIADD[31]) );
    zao211b U1734 ( .A(DW6[0]), .B(QH_PARSE_GO), .C(n2761), .D(n2762), .Y(
        PING_ERR783) );
    zao211b U1735 ( .A(DW7[31]), .B(n2763), .C(n2764), .D(n2765), .Y(TRAN_CMD
        [103]) );
    zao211b U1736 ( .A(DW7[30]), .B(n2763), .C(n2766), .D(n2767), .Y(TRAN_CMD
        [102]) );
    zao211b U1737 ( .A(DW7[29]), .B(n2763), .C(n2768), .D(n2769), .Y(TRAN_CMD
        [101]) );
    zao211b U1738 ( .A(DW7[28]), .B(n2763), .C(n2770), .D(n2771), .Y(TRAN_CMD
        [100]) );
    zao211b U1739 ( .A(n2763), .B(DW7[27]), .C(n2772), .D(n2773), .Y(TRAN_CMD
        [99]) );
    zao211b U1740 ( .A(DW7[26]), .B(n2763), .C(n2774), .D(n2775), .Y(TRAN_CMD
        [98]) );
    zao211b U1741 ( .A(DW7[25]), .B(n2763), .C(n2776), .D(n2777), .Y(TRAN_CMD
        [97]) );
    zao211b U1742 ( .A(DW7[24]), .B(n2763), .C(n2778), .D(n2779), .Y(TRAN_CMD
        [96]) );
    zao211b U1743 ( .A(DW7[23]), .B(n2763), .C(n2780), .D(n2781), .Y(TRAN_CMD
        [95]) );
    zao211b U1744 ( .A(DW7[22]), .B(n2763), .C(n2782), .D(n2783), .Y(TRAN_CMD
        [94]) );
    zao211b U1745 ( .A(DW7[21]), .B(n2763), .C(n2784), .D(n2785), .Y(TRAN_CMD
        [93]) );
    zao211b U1746 ( .A(DW7[20]), .B(n2763), .C(n2786), .D(n2787), .Y(TRAN_CMD
        [92]) );
    zao211b U1747 ( .A(DW7[19]), .B(n2763), .C(n2788), .D(n2789), .Y(TRAN_CMD
        [91]) );
    zao211b U1748 ( .A(DW7[18]), .B(n2763), .C(n2790), .D(n2791), .Y(TRAN_CMD
        [90]) );
    zao211b U1749 ( .A(DW7[17]), .B(n2763), .C(n2792), .D(n2793), .Y(TRAN_CMD
        [89]) );
    zao211b U1750 ( .A(DW7[16]), .B(n2763), .C(n2794), .D(n2795), .Y(TRAN_CMD
        [88]) );
    zao211b U1751 ( .A(DW7[15]), .B(n2763), .C(n2796), .D(n2797), .Y(TRAN_CMD
        [87]) );
    zao211b U1752 ( .A(DW7[14]), .B(n2763), .C(n2798), .D(n2799), .Y(TRAN_CMD
        [86]) );
    zao211b U1753 ( .A(DW7[13]), .B(n2763), .C(n2800), .D(n2801), .Y(TRAN_CMD
        [85]) );
    zao211b U1754 ( .A(DW7[12]), .B(n2763), .C(n2802), .D(n2803), .Y(TRAN_CMD
        [84]) );
    zan4b U1755 ( .A(QHSM[2]), .B(n2888), .C(n2889), .D(n2498), .Y(n2495) );
    zoa21d U1756 ( .A(QHSM[9]), .B(QHSM[6]), .C(PHASENXT_resultwb), .Y(n2893)
         );
    zoa21d U1757 ( .A(UP_DW6[8]), .B(TRAN_CMD[5]), .C(n2515), .Y(n2894) );
    zoa21d U1758 ( .A(n2899), .B(n2900), .C(n2901), .Y(n2898) );
    zoa21d U1759 ( .A(n2907), .B(n2910), .C(n2911), .Y(n2909) );
    zoa21d U1760 ( .A(QHSM[11]), .B(n2921), .C(QHSM[10]), .Y(n2920) );
    zoa21d U1761 ( .A(n2926), .B(n2927), .C(QHSM[2]), .Y(n2925) );
    zoa21d U1762 ( .A(QHSM[0]), .B(QHSM[3]), .C(QHSM[4]), .Y(n2928) );
    zoa21d U1763 ( .A(IMMEDRETRY), .B(n2930), .C(n2931), .Y(n2929) );
    zoa21d U1764 ( .A(RXSTALL), .B(BABBLE), .C(n2521), .Y(n2932) );
    zoa21d U1765 ( .A(n2287), .B(QHSM[5]), .C(n2935), .Y(n2507) );
    zoa21d U1766 ( .A(PARSEQHEND), .B(n2534), .C(n2942), .Y(n2506) );
    zinr2b U1767 ( .A(NAKCNTSM[0]), .B(NAKCNTSM[1]), .Y(n2944) );
    zinr2b U1768 ( .A(NAKCNTSMNXT[0]), .B(NAKCNTSMNXT[1]), .Y(n2945) );
    zoa21d U1769 ( .A(n2949), .B(n2950), .C(n2534), .Y(n2656) );
    zoa21d U1770 ( .A(CACHE_INVALID), .B(n2534), .C(n2942), .Y(n2513) );
    zoa21d U1771 ( .A(SPD), .B(n2957), .C(n2521), .Y(n2956) );
    zoa21d U1772 ( .A(n2299), .B(RXSTALL), .C(n2521), .Y(n2960) );
    zan4b U1773 ( .A(n2511), .B(n2961), .C(ACCEPT_DATA), .D(n2962), .Y(n2957)
         );
    zor3b U1774 ( .A(QHSM[10]), .B(QHSM[11]), .C(n2921), .Y(n2965) );
    zor3b U1775 ( .A(QHSM[4]), .B(QHSM[3]), .C(QHSM[0]), .Y(n2927) );
    zor3b U1776 ( .A(QHSM[4]), .B(QHSM[2]), .C(n2926), .Y(n2968) );
    zor3b U1777 ( .A(QHSM[3]), .B(n2650), .C(n2968), .Y(n2969) );
    zor6b U1778 ( .A(QHSM[10]), .B(CACHEPHASE), .C(n2964), .D(n2970), .E(n2927
        ), .F(QHCIREQ), .Y(n2971) );
    zor3b U1779 ( .A(QHSM[2]), .B(QHSM[1]), .C(n2927), .Y(n2972) );
    zor4b U1780 ( .A(QHSM[5]), .B(n2974), .C(n2508), .D(n2973), .Y(n2916) );
    zor3b U1781 ( .A(QHSM[9]), .B(n2927), .C(n2964), .Y(n2976) );
    zor4b U1782 ( .A(CACHEPHASE), .B(n2977), .C(n2976), .D(QHCIREQ), .Y(n2892)
         );
    zor3b U1783 ( .A(n2971), .B(QRXERR), .C(BABBLE), .Y(n2891) );
    zor3b U1784 ( .A(DW6[9]), .B(UP_DW6[8]), .C(TRAN_CMD[6]), .Y(n2943) );
    zor3b U1785 ( .A(n2328), .B(n3014), .C(n3016), .Y(n3020) );
    zor3b U1786 ( .A(CPAGE_0), .B(n2328), .C(n3014), .Y(n2808) );
    zor3b U1787 ( .A(CPAGE_1), .B(n2328), .C(n3016), .Y(n2806) );
    zor4b U1788 ( .A(BABBLE), .B(n3025), .C(n2903), .D(n2660), .Y(n3024) );
    zor4b U1789 ( .A(QHSM[7]), .B(n3047), .C(n2963), .D(n2973), .Y(n2913) );
    zor4b U1790 ( .A(QHSM[8]), .B(n3048), .C(n2963), .D(n2973), .Y(n2914) );
    zor4b U1791 ( .A(UP_DW5[4]), .B(UP_DW5[3]), .C(UP_DW5[2]), .D(UP_DW5[1]), 
        .Y(n3050) );
    zor5b U1792 ( .A(QHSM[0]), .B(QHSM[3]), .C(QHSM[2]), .D(n3053), .E(n2926), 
        .Y(n3054) );
    zor4b U1793 ( .A(QHSM[6]), .B(n3055), .C(n2508), .D(n2973), .Y(n2917) );
    zor4b U1794 ( .A(QHSM[10]), .B(QHSM[1]), .C(CACHEPHASE), .D(n2976), .Y(
        n3058) );
    zor3b U1795 ( .A(n2325), .B(n2932), .C(n2299), .Y(n2527) );
    zor3b U1796 ( .A(DWCNT[1]), .B(DWCNT[2]), .C(n3066), .Y(n3067) );
    zor3b U1797 ( .A(DWCNT[0]), .B(DWCNT[1]), .C(DWCNT[2]), .Y(n3072) );
    zor3b U1798 ( .A(n3074), .B(n3070), .C(n3066), .Y(n3076) );
    zor3b U1799 ( .A(n3074), .B(n3070), .C(n3069), .Y(n3077) );
    zor3b U1800 ( .A(DWCNT[1]), .B(n3070), .C(n3066), .Y(n3078) );
    zor3b U1801 ( .A(DWCNT[2]), .B(n3074), .C(n3069), .Y(n3079) );
    zor2d U1802 ( .A(n2940), .B(QH_PARSE_GO), .Y(n2662) );
    zor4b U1803 ( .A(n2946), .B(n2940), .C(n2948), .D(n3030), .Y(n2652) );
    zor4b U1804 ( .A(n3083), .B(n3084), .C(n3085), .D(n2899), .Y(n3082) );
    zor2d U1805 ( .A(n3087), .B(n3088), .Y(n2542) );
    zor2d U1806 ( .A(n3061), .B(n3088), .Y(n2540) );
    zor3b U1807 ( .A(n2967), .B(n2650), .C(n2534), .Y(n2504) );
    zao211b U1808 ( .A(BABBLE), .B(n2521), .C(QTDHALT), .D(n2960), .Y(n3096)
         );
    zor3b U1809 ( .A(n2900), .B(n3102), .C(n2299), .Y(n3101) );
    zor4b U1810 ( .A(PIDERR), .B(CRCERR), .C(TMOUT), .D(n2895), .Y(n3108) );
    zao222b U1811 ( .A(DW11[27]), .B(n2327), .C(DW10[27]), .D(n3109), .E(n3110
        ), .F(DW9[27]), .Y(n2773) );
    zao222b U1812 ( .A(DW11[26]), .B(n2327), .C(DW10[26]), .D(n3109), .E(DW9
        [26]), .F(n3110), .Y(n2775) );
    zao222b U1813 ( .A(DW11[25]), .B(n2328), .C(DW10[25]), .D(n3109), .E(DW9
        [25]), .F(n3110), .Y(n2777) );
    zao222b U1814 ( .A(DW11[24]), .B(n2328), .C(DW10[24]), .D(n3109), .E(DW9
        [24]), .F(n3110), .Y(n2779) );
    zao222b U1815 ( .A(DW11[23]), .B(n2327), .C(DW10[23]), .D(n3109), .E(DW9
        [23]), .F(n3110), .Y(n2781) );
    zao222b U1816 ( .A(DW11[22]), .B(n2327), .C(DW10[22]), .D(n3109), .E(DW9
        [22]), .F(n3110), .Y(n2783) );
    zao222b U1817 ( .A(DW11[21]), .B(n2327), .C(DW10[21]), .D(n3109), .E(DW9
        [21]), .F(n3110), .Y(n2785) );
    zao222b U1818 ( .A(DW11[20]), .B(n2327), .C(DW10[20]), .D(n3109), .E(DW9
        [20]), .F(n3110), .Y(n2787) );
    zao222b U1819 ( .A(DW11[19]), .B(n2327), .C(DW10[19]), .D(n3109), .E(DW9
        [19]), .F(n3110), .Y(n2789) );
    zao222b U1820 ( .A(DW11[18]), .B(n2327), .C(DW10[18]), .D(n3109), .E(DW9
        [18]), .F(n3110), .Y(n2791) );
    zao222b U1821 ( .A(DW11[17]), .B(n2328), .C(DW10[17]), .D(n3109), .E(DW9
        [17]), .F(n3110), .Y(n2793) );
    zao222b U1822 ( .A(DW11[16]), .B(n2327), .C(DW10[16]), .D(n3109), .E(DW9
        [16]), .F(n3110), .Y(n2795) );
    zao222b U1823 ( .A(DW11[15]), .B(n2327), .C(DW10[15]), .D(n3109), .E(DW9
        [15]), .F(n3110), .Y(n2797) );
    zao222b U1824 ( .A(DW11[14]), .B(n2327), .C(DW10[14]), .D(n3109), .E(DW9
        [14]), .F(n3110), .Y(n2799) );
    zao222b U1825 ( .A(DW11[13]), .B(n2327), .C(DW10[13]), .D(n3109), .E(DW9
        [13]), .F(n3110), .Y(n2801) );
    zao222b U1826 ( .A(DW11[12]), .B(n2327), .C(DW10[12]), .D(n3109), .E(DW9
        [12]), .F(n3110), .Y(n2803) );
    zao222b U1827 ( .A(DW11[31]), .B(n2327), .C(DW10[31]), .D(n3109), .E(DW9
        [31]), .F(n3110), .Y(n2765) );
    zao222b U1828 ( .A(DW11[30]), .B(n2327), .C(DW10[30]), .D(n3109), .E(DW9
        [30]), .F(n3110), .Y(n2767) );
    zao222b U1829 ( .A(DW11[29]), .B(n2327), .C(DW10[29]), .D(n3109), .E(DW9
        [29]), .F(n3110), .Y(n2769) );
    zao222b U1830 ( .A(DW11[28]), .B(n2327), .C(DW10[28]), .D(n3109), .E(DW9
        [28]), .F(n3110), .Y(n2771) );
    zao222b U1831 ( .A(QHSM[13]), .B(n2358), .C(QHSM[9]), .D(QHCIMWR), .E(QHSM
        [11]), .F(n2921), .Y(n3111) );
    zao211b U1832 ( .A(n3118), .B(n3119), .C(n2928), .D(n2925), .Y(n3117) );
    zao211b U1833 ( .A(PCIEND), .B(n3120), .C(GEN_PERR), .D(n3117), .Y(n2493)
         );
    zao211b U1834 ( .A(TRAN_CMD[7]), .B(n2979), .C(n2959), .D(n3021), .Y(n3102
        ) );
    zao222b U1835 ( .A(DW7[9]), .B(n3172), .C(DW4[9]), .D(n3173), .E(DW3[9]), 
        .F(n3175), .Y(n2692) );
    zao222b U1836 ( .A(DW7[8]), .B(n3123), .C(DW4[8]), .D(n3124), .E(DW3[8]), 
        .F(n3125), .Y(n2689) );
    zao222b U1837 ( .A(DW7[7]), .B(n3171), .C(DW4[7]), .D(n3173), .E(DW3[7]), 
        .F(n3174), .Y(n2686) );
    zao222b U1838 ( .A(DW7[6]), .B(n3172), .C(DW4[6]), .D(n3124), .E(DW3[6]), 
        .F(n3175), .Y(n2683) );
    zao222b U1839 ( .A(DW7[5]), .B(n3123), .C(DW4[5]), .D(n3173), .E(DW3[5]), 
        .F(n3125), .Y(n2680) );
    zao222b U1840 ( .A(DW7[4]), .B(n3171), .C(DW4[4]), .D(n3124), .E(DW3[4]), 
        .F(n3174), .Y(n2677) );
    zao222b U1841 ( .A(DW7[31]), .B(n3172), .C(DW4[31]), .D(n3173), .E(DW3[31]
        ), .F(n3175), .Y(n2758) );
    zao222b U1842 ( .A(DW7[30]), .B(n3123), .C(DW4[30]), .D(n3124), .E(DW3[30]
        ), .F(n3125), .Y(n2755) );
    zao222b U1843 ( .A(DW7[3]), .B(n3171), .C(DW4[3]), .D(n3173), .E(DW3[3]), 
        .F(n3174), .Y(n2674) );
    zao222b U1844 ( .A(DW7[29]), .B(n3172), .C(DW4[29]), .D(n3124), .E(DW3[29]
        ), .F(n3175), .Y(n2752) );
    zao222b U1845 ( .A(DW7[28]), .B(n3123), .C(DW4[28]), .D(n3173), .E(DW3[28]
        ), .F(n3125), .Y(n2749) );
    zao222b U1846 ( .A(DW7[27]), .B(n3171), .C(DW4[27]), .D(n3124), .E(DW3[27]
        ), .F(n3175), .Y(n2746) );
    zao222b U1847 ( .A(DW7[26]), .B(n3172), .C(DW4[26]), .D(n3173), .E(DW3[26]
        ), .F(n3174), .Y(n2743) );
    zao222b U1848 ( .A(DW7[25]), .B(n3123), .C(DW4[25]), .D(n3124), .E(DW3[25]
        ), .F(n3125), .Y(n2740) );
    zao222b U1849 ( .A(DW7[24]), .B(n3172), .C(DW4[24]), .D(n3173), .E(DW3[24]
        ), .F(n3174), .Y(n2737) );
    zao222b U1850 ( .A(DW7[23]), .B(n3123), .C(DW4[23]), .D(n3124), .E(DW3[23]
        ), .F(n3175), .Y(n2734) );
    zao222b U1851 ( .A(DW7[22]), .B(n3171), .C(DW4[22]), .D(n3173), .E(DW3[22]
        ), .F(n3125), .Y(n2731) );
    zao222b U1852 ( .A(DW7[21]), .B(n3171), .C(DW4[21]), .D(n3124), .E(DW3[21]
        ), .F(n3174), .Y(n2728) );
    zao222b U1853 ( .A(DW7[20]), .B(n3172), .C(DW4[20]), .D(n3173), .E(DW3[20]
        ), .F(n3175), .Y(n2725) );
    zao222b U1854 ( .A(DW7[2]), .B(n3123), .C(DW4[2]), .D(n3124), .E(DW3[2]), 
        .F(n3125), .Y(n2671) );
    zao222b U1855 ( .A(DW7[19]), .B(n3171), .C(DW4[19]), .D(n3173), .E(DW3[19]
        ), .F(n3174), .Y(n2722) );
    zao222b U1856 ( .A(DW7[18]), .B(n3172), .C(DW4[18]), .D(n3124), .E(DW3[18]
        ), .F(n3175), .Y(n2719) );
    zao222b U1857 ( .A(DW7[17]), .B(n3123), .C(DW4[17]), .D(n3173), .E(DW3[17]
        ), .F(n3125), .Y(n2716) );
    zao222b U1858 ( .A(DW7[16]), .B(n3171), .C(DW4[16]), .D(n3124), .E(DW3[16]
        ), .F(n3174), .Y(n2713) );
    zao222b U1859 ( .A(DW7[15]), .B(n3172), .C(DW4[15]), .D(n3173), .E(DW3[15]
        ), .F(n3175), .Y(n2710) );
    zao222b U1860 ( .A(DW7[14]), .B(n3123), .C(DW4[14]), .D(n3124), .E(DW3[14]
        ), .F(n3125), .Y(n2707) );
    zao222b U1861 ( .A(DW7[13]), .B(n3172), .C(DW4[13]), .D(n3173), .E(DW3[13]
        ), .F(n3174), .Y(n2704) );
    zao222b U1862 ( .A(DW7[12]), .B(n3123), .C(DW4[12]), .D(n3124), .E(DW3[12]
        ), .F(n3175), .Y(n2701) );
    zao222b U1863 ( .A(DW7[11]), .B(n3171), .C(DW4[11]), .D(n3173), .E(DW3[11]
        ), .F(n3125), .Y(n2698) );
    zao222b U1864 ( .A(DW7[10]), .B(n3171), .C(DW4[10]), .D(n3124), .E(DW3[10]
        ), .F(n3174), .Y(n2695) );
    zao222b U1865 ( .A(DW7[1]), .B(n3172), .C(DW4[1]), .D(n3173), .E(DW3[1]), 
        .F(n3175), .Y(n2668) );
    zao222b U1866 ( .A(DW7[0]), .B(n3123), .C(n3124), .D(DW4[0]), .E(DW3[0]), 
        .F(n3125), .Y(n2665) );
    zor6b U1867 ( .A(MAXLEN[7]), .B(MAXLEN[6]), .C(MAXLEN[5]), .D(MAXLEN[10]), 
        .E(MAXLEN[9]), .F(MAXLEN[8]), .Y(n2934) );
    zoa21d U1868 ( .A(n2944), .B(n2945), .C(n3132), .Y(n2947) );
    zoai22d U1869 ( .A(RXNYET), .B(n3021), .C(n2515), .D(n2510), .Y(n3133) );
    zan4b U1870 ( .A(n3042), .B(n3033), .C(n3031), .D(n3039), .Y(n3134) );
    zan4b U1871 ( .A(n3037), .B(n3036), .C(n3034), .D(n3032), .Y(n3136) );
    zor3b U1872 ( .A(n2980), .B(n2943), .C(TRAN_CMD[5]), .Y(n2906) );
    zor3b U1873 ( .A(QHSM[4]), .B(n3056), .C(TRAN_CMD[5]), .Y(n2659) );
    zor3b U1874 ( .A(n3133), .B(n3044), .C(n2660), .Y(n2953) );
    zivh U1875 ( .A(n3081), .Y(n2655) );
    zao222b U1876 ( .A(FEMPTY), .B(n3146), .C(n3145), .D(n3150), .E(n3144), 
        .F(n2512), .Y(n2978) );
    zao211b U1877 ( .A(TRAN_CMD[7]), .B(n3021), .C(n3025), .D(n2894), .Y(n3151
        ) );
    zao211b U1878 ( .A(RXNYET), .B(n3151), .C(n2897), .D(n3108), .Y(n3022) );
    zor4b U1879 ( .A(n2905), .B(n2896), .C(n2899), .D(n2660), .Y(n2911) );
    zor4b U1880 ( .A(DW1[31]), .B(DW1[30]), .C(DW1[29]), .D(DW1[28]), .Y(n3132
        ) );
    zao222b U1881 ( .A(IMMEDRETRY), .B(n2294), .C(n3143), .D(n2514), .E(n2293), 
        .F(n3154), .Y(n3057) );
    zao222b U1882 ( .A(n2295), .B(n2501), .C(n2294), .D(n3052), .E(
        CACHE_MODIFY), .F(n3155), .Y(n3137) );
    zor4b U1883 ( .A(n2920), .B(n3111), .C(n3112), .D(n3121), .Y(n3119) );
    zor4b U1884 ( .A(n2288), .B(DW6[6]), .C(n2534), .D(n2922), .Y(n2492) );
    zao211b U1885 ( .A(n2295), .B(ACTIVE), .C(n2296), .D(n2924), .Y(n3120) );
    zor4b U1886 ( .A(n3059), .B(ACTIVE), .C(n3062), .D(QHSMNXT_13), .Y(n3064)
         );
    zao32d U1887 ( .A(n2323), .B(n3070), .C(n3147), .D(n3141), .E(QHDWNUM[0]), 
        .Y(n3127) );
    zao22d U1888 ( .A(n3141), .B(QHDWNUM[3]), .C(DWCNT[3]), .D(n3072), .Y(
        n3125) );
    zao32d U1889 ( .A(n2324), .B(n3074), .C(n3149), .D(n3142), .E(QHDWNUM[0]), 
        .Y(n3123) );
    zor4b U1890 ( .A(TDMAEND), .B(n2524), .C(TRAN_CMD[5]), .D(n2933), .Y(n2935
        ) );
    zoai21d U1891 ( .A(ACCEPT_DATA), .B(n2938), .C(n3104), .Y(n2654) );
    zao32d U1892 ( .A(n3140), .B(TRAN_CMD[5]), .C(ACCEPT_DATA), .D(n3104), .E(
        n2899), .Y(n2653) );
    zor3b U1893 ( .A(CPAGE_1), .B(CPAGE_0), .C(n3012), .Y(n3094) );
    zor3b U1894 ( .A(CACHE_MODIFY), .B(QHSM[2]), .C(PHASENXT_resultwb), .Y(
        n2533) );
    zmux21ld U1895 ( .A(n2524), .B(n3025), .S(UP_DW6[8]), .Y(n2661) );
    zor3b U1896 ( .A(n2959), .B(n2314), .C(n2956), .Y(n3107) );
    zor2d U1897 ( .A(n3061), .B(n3088), .Y(n3161) );
    zor2d U1898 ( .A(n3061), .B(n3088), .Y(n3162) );
    zor2d U1899 ( .A(n3087), .B(n3088), .Y(n3163) );
    zor2d U1900 ( .A(n3087), .B(n3088), .Y(n3164) );
    zor3b U1901 ( .A(CPAGE_1), .B(CPAGE_0), .C(n2328), .Y(n3165) );
    zor3b U1902 ( .A(CPAGE_1), .B(n2328), .C(n3016), .Y(n3166) );
    zor3b U1903 ( .A(CPAGE_1), .B(n2328), .C(n3016), .Y(n3167) );
    zor3b U1904 ( .A(CPAGE_0), .B(n2328), .C(n3014), .Y(n3168) );
    zor3b U1905 ( .A(CPAGE_0), .B(n2328), .C(n3014), .Y(n3169) );
    zao32d U1906 ( .A(DWCNT[2]), .B(n3074), .C(n3149), .D(n3142), .E(QHDWNUM
        [0]), .Y(n3171) );
    zao32d U1907 ( .A(n2324), .B(n3074), .C(n3149), .D(n3142), .E(QHDWNUM[0]), 
        .Y(n3172) );
    zao22d U1908 ( .A(n3141), .B(QHDWNUM[3]), .C(DWCNT[3]), .D(n3072), .Y(
        n3174) );
    zao22d U1909 ( .A(n3141), .B(QHDWNUM[3]), .C(DWCNT[3]), .D(n3072), .Y(
        n3175) );
    zao32d U1910 ( .A(DWCNT[1]), .B(n3070), .C(n3147), .D(n3141), .E(QHDWNUM
        [0]), .Y(n3177) );
    zao32d U1911 ( .A(n2323), .B(n3070), .C(n3147), .D(n3141), .E(QHDWNUM[0]), 
        .Y(n3178) );
    zor3b U1912 ( .A(DWCNT[2]), .B(n3074), .C(n3069), .Y(n3179) );
    zor3b U1913 ( .A(DWCNT[2]), .B(n3074), .C(n3069), .Y(n3180) );
    zor3b U1914 ( .A(DWCNT[1]), .B(n3070), .C(n3066), .Y(n3181) );
    zor3b U1915 ( .A(DWCNT[1]), .B(n3070), .C(n3066), .Y(n3182) );
    zor3b U1916 ( .A(n3074), .B(n3070), .C(n3069), .Y(n3183) );
    zor3b U1917 ( .A(n3074), .B(n3070), .C(n3069), .Y(n3184) );
    zor3b U1918 ( .A(n3074), .B(n3070), .C(n3066), .Y(n3185) );
    zor3b U1919 ( .A(n3074), .B(n3070), .C(n3066), .Y(n3186) );
endmodule


module ASYNC_MUX ( QH_CACHE_EN1, QH_CACHE_EN2, DWNUM, QHDWNUM1, QHDWNUM2, 
    EDWNUM, DWOFFSET, QDWOFFSET1, QDWOFFSET2, EDWOFFSET, EHCI_MAC_EOT, 
    QHCIGNT1, QHCIGNT2, QHCIMWR1, QHCIMWR2, HCIMWR, PCIEND, QPCIEND1, QPCIEND2, 
    QH_ACT1, QH_ACT2, QH_MAC_EOT1, QH_MAC_EOT2, USBDMA_SEL, CRCERR, BABBLE, 
    PIDERR, TMOUT, TOGMATCH, RXNAK, RXNYET, RXSTALL, RXACK, RXDATA0, RXDATA1, 
    RXPIDERR, SPD, ACTLEN, CRCERR1, BABBLE1, PIDERR1, TMOUT1, TOGMATCH1, 
    RXNAK1, RXNYET1, RXSTALL1, RXACK1, RXDATA01, RXDATA11, RXPIDERR1, SPD1, 
    ACTLEN1, CRCERR2, BABBLE2, PIDERR2, TMOUT2, TOGMATCH2, RXNAK2, RXNYET2, 
    RXSTALL2, RXACK2, RXDATA02, RXDATA12, RXPIDERR2, SPD2, ACTLEN2 );
input  [3:0] DWNUM;
input  [3:0] QHDWNUM1;
input  [3:0] DWOFFSET;
output [10:0] ACTLEN1;
input  [4:0] USBDMA_SEL;
input  [3:0] QHDWNUM2;
output [3:0] EDWNUM;
input  [3:0] QDWOFFSET1;
output [3:0] EDWOFFSET;
input  [10:0] ACTLEN;
output [10:0] ACTLEN2;
input  [3:0] QDWOFFSET2;
input  QH_CACHE_EN1, QH_CACHE_EN2, EHCI_MAC_EOT, QHCIGNT1, QHCIGNT2, QHCIMWR1, 
    QHCIMWR2, PCIEND, QH_ACT1, QH_ACT2, CRCERR, BABBLE, PIDERR, TMOUT, 
    TOGMATCH, RXNAK, RXNYET, RXSTALL, RXACK, RXDATA0, RXDATA1, RXPIDERR, SPD;
output HCIMWR, QPCIEND1, QPCIEND2, QH_MAC_EOT1, QH_MAC_EOT2, CRCERR1, BABBLE1, 
    PIDERR1, TMOUT1, TOGMATCH1, RXNAK1, RXNYET1, RXSTALL1, RXACK1, RXDATA01, 
    RXDATA11, RXPIDERR1, SPD1, CRCERR2, BABBLE2, PIDERR2, TMOUT2, TOGMATCH2, 
    RXNAK2, RXNYET2, RXSTALL2, RXACK2, RXDATA02, RXDATA12, RXPIDERR2, SPD2;
    wire n723, n724, n725;
    zan2b U39 ( .A(CRCERR), .B(USBDMA_SEL[3]), .Y(CRCERR2) );
    zan2b U40 ( .A(BABBLE), .B(USBDMA_SEL[3]), .Y(BABBLE2) );
    zan2b U41 ( .A(PIDERR), .B(USBDMA_SEL[3]), .Y(PIDERR2) );
    zan2b U42 ( .A(TMOUT), .B(USBDMA_SEL[3]), .Y(TMOUT2) );
    zan2b U43 ( .A(USBDMA_SEL[3]), .B(TOGMATCH), .Y(TOGMATCH2) );
    zan2b U44 ( .A(RXNAK), .B(USBDMA_SEL[3]), .Y(RXNAK2) );
    zan2b U45 ( .A(RXNYET), .B(USBDMA_SEL[3]), .Y(RXNYET2) );
    zan2b U46 ( .A(RXSTALL), .B(USBDMA_SEL[3]), .Y(RXSTALL2) );
    zan2b U47 ( .A(RXACK), .B(USBDMA_SEL[3]), .Y(RXACK2) );
    zan2b U48 ( .A(RXDATA0), .B(USBDMA_SEL[3]), .Y(RXDATA02) );
    zan2b U49 ( .A(RXDATA1), .B(USBDMA_SEL[3]), .Y(RXDATA12) );
    zan2b U50 ( .A(RXPIDERR), .B(USBDMA_SEL[3]), .Y(RXPIDERR2) );
    zan2b U51 ( .A(SPD), .B(USBDMA_SEL[3]), .Y(SPD2) );
    zan2b U52 ( .A(ACTLEN[10]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[10]) );
    zan2b U53 ( .A(ACTLEN[9]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[9]) );
    zan2b U54 ( .A(ACTLEN[8]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[8]) );
    zan2b U55 ( .A(ACTLEN[7]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[7]) );
    zan2b U56 ( .A(ACTLEN[6]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[6]) );
    zan2b U57 ( .A(ACTLEN[5]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[5]) );
    zan2b U58 ( .A(ACTLEN[4]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[4]) );
    zan2b U59 ( .A(ACTLEN[3]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[3]) );
    zan2b U60 ( .A(ACTLEN[2]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[2]) );
    zan2b U61 ( .A(ACTLEN[1]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[1]) );
    zan2b U62 ( .A(ACTLEN[0]), .B(USBDMA_SEL[3]), .Y(ACTLEN2[0]) );
    zao222b U63 ( .A(QDWOFFSET2[3]), .B(n723), .C(DWOFFSET[3]), .D(n724), .E(
        QH_CACHE_EN1), .F(QDWOFFSET1[3]), .Y(EDWOFFSET[3]) );
    zao222b U64 ( .A(QDWOFFSET2[2]), .B(n723), .C(DWOFFSET[2]), .D(n724), .E(
        QDWOFFSET1[2]), .F(QH_CACHE_EN1), .Y(EDWOFFSET[2]) );
    zao222b U65 ( .A(QDWOFFSET2[1]), .B(n723), .C(DWOFFSET[1]), .D(n724), .E(
        QDWOFFSET1[1]), .F(QH_CACHE_EN1), .Y(EDWOFFSET[1]) );
    zao222b U66 ( .A(QDWOFFSET2[0]), .B(n723), .C(DWOFFSET[0]), .D(n724), .E(
        QDWOFFSET1[0]), .F(QH_CACHE_EN1), .Y(EDWOFFSET[0]) );
    zan2b U67 ( .A(CRCERR), .B(USBDMA_SEL[2]), .Y(CRCERR1) );
    zan2b U68 ( .A(BABBLE), .B(USBDMA_SEL[2]), .Y(BABBLE1) );
    zan2b U69 ( .A(PIDERR), .B(USBDMA_SEL[2]), .Y(PIDERR1) );
    zan2b U70 ( .A(TMOUT), .B(USBDMA_SEL[2]), .Y(TMOUT1) );
    zan2b U71 ( .A(USBDMA_SEL[2]), .B(TOGMATCH), .Y(TOGMATCH1) );
    zan2b U72 ( .A(RXNAK), .B(USBDMA_SEL[2]), .Y(RXNAK1) );
    zan2b U73 ( .A(RXNYET), .B(USBDMA_SEL[2]), .Y(RXNYET1) );
    zan2b U74 ( .A(RXSTALL), .B(USBDMA_SEL[2]), .Y(RXSTALL1) );
    zan2b U75 ( .A(RXACK), .B(USBDMA_SEL[2]), .Y(RXACK1) );
    zan2b U76 ( .A(RXDATA0), .B(USBDMA_SEL[2]), .Y(RXDATA01) );
    zan2b U77 ( .A(RXDATA1), .B(USBDMA_SEL[2]), .Y(RXDATA11) );
    zan2b U78 ( .A(RXPIDERR), .B(USBDMA_SEL[2]), .Y(RXPIDERR1) );
    zan2b U79 ( .A(SPD), .B(USBDMA_SEL[2]), .Y(SPD1) );
    zan2b U80 ( .A(ACTLEN[10]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[10]) );
    zan2b U81 ( .A(ACTLEN[9]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[9]) );
    zan2b U82 ( .A(ACTLEN[8]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[8]) );
    zan2b U83 ( .A(ACTLEN[7]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[7]) );
    zan2b U84 ( .A(ACTLEN[6]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[6]) );
    zan2b U85 ( .A(ACTLEN[5]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[5]) );
    zan2b U86 ( .A(ACTLEN[4]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[4]) );
    zan2b U87 ( .A(ACTLEN[3]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[3]) );
    zan2b U88 ( .A(ACTLEN[2]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[2]) );
    zan2b U89 ( .A(ACTLEN[1]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[1]) );
    zan2b U90 ( .A(ACTLEN[0]), .B(USBDMA_SEL[2]), .Y(ACTLEN1[0]) );
    zao222b U91 ( .A(QHDWNUM2[3]), .B(QHCIGNT2), .C(DWNUM[3]), .D(n725), .E(
        QHDWNUM1[3]), .F(QHCIGNT1), .Y(EDWNUM[3]) );
    zao222b U92 ( .A(QHDWNUM1[0]), .B(QHCIGNT1), .C(DWNUM[0]), .D(n725), .E(
        QHDWNUM2[0]), .F(QHCIGNT2), .Y(EDWNUM[0]) );
    zan2b U93 ( .A(QH_ACT1), .B(EHCI_MAC_EOT), .Y(QH_MAC_EOT1) );
    zan2b U94 ( .A(EHCI_MAC_EOT), .B(QH_ACT2), .Y(QH_MAC_EOT2) );
    zao222b U95 ( .A(QHDWNUM1[1]), .B(QHCIGNT1), .C(DWNUM[1]), .D(n725), .E(
        QHDWNUM2[1]), .F(QHCIGNT2), .Y(EDWNUM[1]) );
    zan2b U96 ( .A(QHCIGNT1), .B(PCIEND), .Y(QPCIEND1) );
    zao222b U97 ( .A(QHDWNUM2[2]), .B(QHCIGNT2), .C(DWNUM[2]), .D(n725), .E(
        QHDWNUM1[2]), .F(QHCIGNT1), .Y(EDWNUM[2]) );
    zan2b U98 ( .A(QHCIGNT2), .B(PCIEND), .Y(QPCIEND2) );
    zao22b U99 ( .A(QHCIMWR1), .B(QHCIGNT1), .C(QHCIMWR2), .D(QHCIGNT2), .Y(
        HCIMWR) );
    znr2b U100 ( .A(QH_CACHE_EN2), .B(QH_CACHE_EN1), .Y(n724) );
    zinr2b U101 ( .A(QH_CACHE_EN2), .B(QH_CACHE_EN1), .Y(n723) );
    znr2b U102 ( .A(QHCIGNT2), .B(QHCIGNT1), .Y(n725) );
endmodule


module ASYNC_ADCTL ( PCICLK, TRST_, DWCNT, WR_ASYNCADDR, RUN, ADI, ASYNC_ACT, 
    ASYNC_EN, ASYNCLISTADDR, DW1_0, DW2_0, PARSEQHEND1, PARSEQHEND2, QHCIGNT1, 
    QHCIGNT2, QHCIADR1, QHCIADR2, HCIADR, QHCIADD1, QHCIADD2, HCIADD, 
    ASYNC_EMPTY1, ASYNC_EMPTY2 );
input  [3:0] DWCNT;
input  [31:0] ADI;
input  [31:0] QHCIADD1;
input  [31:0] DW2_0;
input  [31:0] QHCIADR1;
output [31:0] ASYNCLISTADDR;
input  [31:0] DW1_0;
input  [31:0] QHCIADR2;
output [31:0] HCIADR;
input  [31:0] QHCIADD2;
output [31:0] HCIADD;
input  PCICLK, TRST_, WR_ASYNCADDR, RUN, ASYNC_ACT, ASYNC_EN, PARSEQHEND1, 
    PARSEQHEND2, QHCIGNT1, QHCIGNT2, ASYNC_EMPTY1, ASYNC_EMPTY2;
    wire ASYNCLISTADDR136_15, SPAREO6, HCIADR_p_2, ASYNCLISTADDR136_29, 
        HCIADR_p_13, ASYNCLISTADDR136_3, HCIADR_p_26, ASYNCLISTADDR136_20, 
        ASYNCLISTADDR136_27, SPAREO0_, SPAREO8, HCIADR_p_21, HCIADR_p_14, 
        ASYNCLISTADDR136_4, HCIADR_p_5, SPAREO1, HCIADR_p_28, 
        ASYNCLISTADDR136_12, HCIADR_p_20, SPAREO9, ASYNCLISTADDR136_26, 
        HCIADR_p_29, ASYNCLISTADDR136_13, SPAREO0, HCIADR_p_4, HCIADR_p_15, 
        ASYNCLISTADDR136_5, ASYNCLISTADDR136_28, HCIADR_p_12, 
        ASYNCLISTADDR136_2, HCIADR_p_3, SPAREO7, ASYNCLISTADDR136_14, 
        ASYNCLISTADDR136_21, HCIADR_p_27, ASYNCLISTADDR136_31, 
        ASYNCLISTADDR136_16, SPAREO5, HCIADR_p_1, ASYNCLISTADDR136_0, 
        HCIADR_p_10, HCIADR_p_25, HCIADR_p_8, ASYNCLISTADDR136_9, 
        ASYNCLISTADDR136_23, HCIADR_p_19, ASYNCLISTADDR136_24, HCIADR_p_22, 
        ASYNCLISTADDR136_18, ASYNCLISTADDR136_7, HCIADR_p_17, HCIADR_p_6, 
        SPAREO2, ASYNCLISTADDR136_11, HCIADR_p_23, ASYNCLISTADDR136_19, 
        ASYNCLISTADDR136_25, ASYNCLISTADDR136_10, SPAREO3, SPAREO1_, 
        HCIADR_p_7, ASYNCLISTADDR136_6, HCIADR_p_16, ASYNCLISTADDR136_1, 
        HCIADR_p_11, HCIADR_p_0, SPAREO4, ASYNCLISTADDR136_30, 
        ASYNCLISTADDR136_17, ASYNCLISTADDR136_8, ASYNCLISTADDR136_22, 
        HCIADR_p_18, ASYNCADDR_WE, HCIADR_p_9, HCIADR_p_24, n241, n242, n243, 
        n244, n245, n246, n247, n248, add_50_carry_29, add_50_carry_1, 
        add_50_carry_20, add_50_carry_15, add_50_carry_8, add_50_carry_28, 
        add_50_carry_27, add_50_carry_26, add_50_carry_12, add_50_carry_6, 
        add_50_carry_14, add_50_carry_13, add_50_carry_7, add_50_carry_24, 
        add_50_carry_23, add_50_carry_21, add_50_carry_16, add_50_carry_9, 
        add_50_carry_2, add_50_carry_18, add_50_carry_25, add_50_carry_11, 
        add_50_carry_5, add_50_carry_19, add_50_carry_10, add_50_carry_4, 
        add_50_carry_22, add_50_carry_17, add_50_carry_3, n249, n250, n251, 
        n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
        n264, n265, n266, n267, n268, n269, n270;
    assign HCIADR[1] = 1'b0;
    assign HCIADR[0] = 1'b0;
    zivb SPARE857 ( .A(SPAREO4), .Y(SPAREO5) );
    znd3b SPARE859 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE850 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE858 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE851 ( .CK(PCICLK), .D(SPAREO7), .R(TRST_), .Q(SPAREO1), .QN(
        SPAREO1_) );
    znr3b SPARE856 ( .A(SPAREO2), .B(ASYNCADDR_WE), .C(SPAREO0_), .Y(SPAREO4)
         );
    zoai21b SPARE854 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE853 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zaoi211b SPARE852 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE855 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zor2b U82 ( .A(n268), .B(n244), .Y(n258) );
    zivc U83 ( .A(n263), .Y(n251) );
    zivc U84 ( .A(n263), .Y(ASYNCADDR_WE) );
    zivb U85 ( .A(n257), .Y(n261) );
    zivb U86 ( .A(PARSEQHEND2), .Y(n256) );
    zan2b U87 ( .A(n250), .B(ASYNCLISTADDR[4]), .Y(ASYNCLISTADDR136_4) );
    zan2b U88 ( .A(n265), .B(ASYNCLISTADDR[3]), .Y(ASYNCLISTADDR136_3) );
    zan2b U89 ( .A(n265), .B(ASYNCLISTADDR[2]), .Y(ASYNCLISTADDR136_2) );
    zan2b U90 ( .A(ASYNCLISTADDR[1]), .B(n265), .Y(ASYNCLISTADDR136_1) );
    zan2b U91 ( .A(ASYNCLISTADDR[0]), .B(n250), .Y(ASYNCLISTADDR136_0) );
    zivc U92 ( .A(n264), .Y(n250) );
    zoai21b U93 ( .A(n255), .B(n259), .C(n263), .Y(n264) );
    zivb U94 ( .A(ASYNC_ACT), .Y(n259) );
    zivc U95 ( .A(n264), .Y(n265) );
    zao22b U96 ( .A(QHCIADD2[1]), .B(n245), .C(QHCIADD1[1]), .D(n268), .Y(
        HCIADD[1]) );
    zao22b U97 ( .A(QHCIADD2[9]), .B(n245), .C(QHCIADD1[9]), .D(n268), .Y(
        HCIADD[9]) );
    zao22b U98 ( .A(QHCIADD1[12]), .B(n246), .C(QHCIADD2[12]), .D(n245), .Y(
        HCIADD[12]) );
    zao22b U99 ( .A(QHCIADD2[14]), .B(n245), .C(QHCIADD1[14]), .D(n246), .Y(
        HCIADD[14]) );
    zao22b U100 ( .A(QHCIADD2[16]), .B(n244), .C(QHCIADD1[16]), .D(n268), .Y(
        HCIADD[16]) );
    zao22b U101 ( .A(QHCIADD2[17]), .B(n244), .C(QHCIADD1[17]), .D(n268), .Y(
        HCIADD[17]) );
    zao22b U102 ( .A(QHCIADD2[21]), .B(n266), .C(QHCIADD1[21]), .D(n268), .Y(
        HCIADD[21]) );
    zao22b U103 ( .A(QHCIADD2[28]), .B(n266), .C(QHCIADD1[28]), .D(n268), .Y(
        HCIADD[28]) );
    zao22b U104 ( .A(QHCIADD2[29]), .B(n244), .C(QHCIADD1[29]), .D(n268), .Y(
        HCIADD[29]) );
    zivc U105 ( .A(n241), .Y(n268) );
    zao22b U106 ( .A(QHCIADD1[31]), .B(n246), .C(QHCIADD2[31]), .D(n266), .Y(
        HCIADD[31]) );
    zivc U107 ( .A(n243), .Y(n267) );
    zivc U108 ( .A(n258), .Y(n249) );
    zivc U109 ( .A(n258), .Y(n270) );
    zdffqrb ASYNCLISTADDR_reg_31 ( .CK(PCICLK), .D(ASYNCLISTADDR136_31), .R(
        TRST_), .Q(ASYNCLISTADDR[31]) );
    zdffqrb ASYNCLISTADDR_reg_30 ( .CK(PCICLK), .D(ASYNCLISTADDR136_30), .R(
        TRST_), .Q(ASYNCLISTADDR[30]) );
    zdffqrb ASYNCLISTADDR_reg_29 ( .CK(PCICLK), .D(ASYNCLISTADDR136_29), .R(
        TRST_), .Q(ASYNCLISTADDR[29]) );
    zdffqrb ASYNCLISTADDR_reg_28 ( .CK(PCICLK), .D(ASYNCLISTADDR136_28), .R(
        TRST_), .Q(ASYNCLISTADDR[28]) );
    zdffqrb ASYNCLISTADDR_reg_27 ( .CK(PCICLK), .D(ASYNCLISTADDR136_27), .R(
        TRST_), .Q(ASYNCLISTADDR[27]) );
    zdffqrb ASYNCLISTADDR_reg_26 ( .CK(PCICLK), .D(ASYNCLISTADDR136_26), .R(
        TRST_), .Q(ASYNCLISTADDR[26]) );
    zdffqrb ASYNCLISTADDR_reg_25 ( .CK(PCICLK), .D(ASYNCLISTADDR136_25), .R(
        TRST_), .Q(ASYNCLISTADDR[25]) );
    zdffqrb ASYNCLISTADDR_reg_24 ( .CK(PCICLK), .D(ASYNCLISTADDR136_24), .R(
        TRST_), .Q(ASYNCLISTADDR[24]) );
    zdffqrb ASYNCLISTADDR_reg_23 ( .CK(PCICLK), .D(ASYNCLISTADDR136_23), .R(
        TRST_), .Q(ASYNCLISTADDR[23]) );
    zdffqrb ASYNCLISTADDR_reg_22 ( .CK(PCICLK), .D(ASYNCLISTADDR136_22), .R(
        TRST_), .Q(ASYNCLISTADDR[22]) );
    zdffqrb ASYNCLISTADDR_reg_21 ( .CK(PCICLK), .D(ASYNCLISTADDR136_21), .R(
        TRST_), .Q(ASYNCLISTADDR[21]) );
    zdffqrb ASYNCLISTADDR_reg_20 ( .CK(PCICLK), .D(ASYNCLISTADDR136_20), .R(
        TRST_), .Q(ASYNCLISTADDR[20]) );
    zdffqrb ASYNCLISTADDR_reg_19 ( .CK(PCICLK), .D(ASYNCLISTADDR136_19), .R(
        TRST_), .Q(ASYNCLISTADDR[19]) );
    zdffqrb ASYNCLISTADDR_reg_18 ( .CK(PCICLK), .D(ASYNCLISTADDR136_18), .R(
        TRST_), .Q(ASYNCLISTADDR[18]) );
    zdffqrb ASYNCLISTADDR_reg_17 ( .CK(PCICLK), .D(ASYNCLISTADDR136_17), .R(
        TRST_), .Q(ASYNCLISTADDR[17]) );
    zdffqrb ASYNCLISTADDR_reg_16 ( .CK(PCICLK), .D(ASYNCLISTADDR136_16), .R(
        TRST_), .Q(ASYNCLISTADDR[16]) );
    zdffqrb ASYNCLISTADDR_reg_15 ( .CK(PCICLK), .D(ASYNCLISTADDR136_15), .R(
        TRST_), .Q(ASYNCLISTADDR[15]) );
    zdffqrb ASYNCLISTADDR_reg_14 ( .CK(PCICLK), .D(ASYNCLISTADDR136_14), .R(
        TRST_), .Q(ASYNCLISTADDR[14]) );
    zdffqrb ASYNCLISTADDR_reg_13 ( .CK(PCICLK), .D(ASYNCLISTADDR136_13), .R(
        TRST_), .Q(ASYNCLISTADDR[13]) );
    zdffqrb ASYNCLISTADDR_reg_12 ( .CK(PCICLK), .D(ASYNCLISTADDR136_12), .R(
        TRST_), .Q(ASYNCLISTADDR[12]) );
    zdffqrb ASYNCLISTADDR_reg_11 ( .CK(PCICLK), .D(ASYNCLISTADDR136_11), .R(
        TRST_), .Q(ASYNCLISTADDR[11]) );
    zdffqrb ASYNCLISTADDR_reg_10 ( .CK(PCICLK), .D(ASYNCLISTADDR136_10), .R(
        TRST_), .Q(ASYNCLISTADDR[10]) );
    zdffqrb ASYNCLISTADDR_reg_9 ( .CK(PCICLK), .D(ASYNCLISTADDR136_9), .R(
        TRST_), .Q(ASYNCLISTADDR[9]) );
    zdffqrb ASYNCLISTADDR_reg_8 ( .CK(PCICLK), .D(ASYNCLISTADDR136_8), .R(
        TRST_), .Q(ASYNCLISTADDR[8]) );
    zdffqrb ASYNCLISTADDR_reg_7 ( .CK(PCICLK), .D(ASYNCLISTADDR136_7), .R(
        TRST_), .Q(ASYNCLISTADDR[7]) );
    zdffqrb ASYNCLISTADDR_reg_6 ( .CK(PCICLK), .D(ASYNCLISTADDR136_6), .R(
        TRST_), .Q(ASYNCLISTADDR[6]) );
    zdffqrb ASYNCLISTADDR_reg_5 ( .CK(PCICLK), .D(ASYNCLISTADDR136_5), .R(
        TRST_), .Q(ASYNCLISTADDR[5]) );
    zdffqrb ASYNCLISTADDR_reg_4 ( .CK(PCICLK), .D(ASYNCLISTADDR136_4), .R(
        TRST_), .Q(ASYNCLISTADDR[4]) );
    zdffqrb ASYNCLISTADDR_reg_3 ( .CK(PCICLK), .D(ASYNCLISTADDR136_3), .R(
        TRST_), .Q(ASYNCLISTADDR[3]) );
    zdffqrb ASYNCLISTADDR_reg_2 ( .CK(PCICLK), .D(ASYNCLISTADDR136_2), .R(
        TRST_), .Q(ASYNCLISTADDR[2]) );
    zdffqrb ASYNCLISTADDR_reg_1 ( .CK(PCICLK), .D(ASYNCLISTADDR136_1), .R(
        TRST_), .Q(ASYNCLISTADDR[1]) );
    zdffqrb ASYNCLISTADDR_reg_0 ( .CK(PCICLK), .D(ASYNCLISTADDR136_0), .R(
        TRST_), .Q(ASYNCLISTADDR[0]) );
    ziv11d U110 ( .A(QHCIGNT1), .Y(n241), .Z(n242) );
    ziv11d U111 ( .A(QHCIGNT2), .Y(n243), .Z(n244) );
    zivc U112 ( .A(n243), .Y(n245) );
    zao22b U113 ( .A(QHCIADD2[0]), .B(n266), .C(QHCIADD1[0]), .D(n268), .Y(
        HCIADD[0]) );
    zao22b U114 ( .A(QHCIADD2[22]), .B(n244), .C(QHCIADD1[22]), .D(n242), .Y(
        HCIADD[22]) );
    zao22b U115 ( .A(QHCIADD2[23]), .B(n266), .C(QHCIADD1[23]), .D(n268), .Y(
        HCIADD[23]) );
    zao22b U116 ( .A(QHCIADD2[4]), .B(n245), .C(QHCIADD1[4]), .D(n268), .Y(
        HCIADD[4]) );
    zao22b U117 ( .A(QHCIADD2[20]), .B(n244), .C(QHCIADD1[20]), .D(n268), .Y(
        HCIADD[20]) );
    zao22b U118 ( .A(QHCIADD2[2]), .B(n266), .C(QHCIADD1[2]), .D(n268), .Y(
        HCIADD[2]) );
    zao22b U119 ( .A(QHCIADD2[15]), .B(n245), .C(QHCIADD1[15]), .D(n268), .Y(
        HCIADD[15]) );
    zao22b U120 ( .A(QHCIADD2[7]), .B(n244), .C(QHCIADD1[7]), .D(n268), .Y(
        HCIADD[7]) );
    zao22b U121 ( .A(QHCIADD1[19]), .B(n269), .C(QHCIADD2[19]), .D(n245), .Y(
        HCIADD[19]) );
    zao22b U122 ( .A(QHCIADD1[6]), .B(n242), .C(QHCIADD2[6]), .D(n266), .Y(
        HCIADD[6]) );
    zao22b U123 ( .A(QHCIADD1[24]), .B(n242), .C(QHCIADD2[24]), .D(n244), .Y(
        HCIADD[24]) );
    zao22b U124 ( .A(QHCIADD1[3]), .B(n269), .C(QHCIADD2[3]), .D(n244), .Y(
        HCIADD[3]) );
    zao22b U125 ( .A(QHCIADD1[18]), .B(n246), .C(QHCIADD2[18]), .D(n266), .Y(
        HCIADD[18]) );
    zao22b U126 ( .A(QHCIADD1[26]), .B(n269), .C(QHCIADD2[26]), .D(n245), .Y(
        HCIADD[26]) );
    zao22b U127 ( .A(QHCIADD1[11]), .B(n242), .C(QHCIADD2[11]), .D(n245), .Y(
        HCIADD[11]) );
    zao22b U128 ( .A(QHCIADD1[8]), .B(n269), .C(QHCIADD2[8]), .D(n266), .Y(
        HCIADD[8]) );
    zivc U129 ( .A(n243), .Y(n266) );
    zivc U130 ( .A(n241), .Y(n246) );
    zao22b U131 ( .A(QHCIADD1[30]), .B(n246), .C(QHCIADD2[30]), .D(n266), .Y(
        HCIADD[30]) );
    zao22b U132 ( .A(QHCIADD1[13]), .B(n269), .C(QHCIADD2[13]), .D(n244), .Y(
        HCIADD[13]) );
    zao22b U133 ( .A(QHCIADD1[27]), .B(n269), .C(QHCIADD2[27]), .D(n244), .Y(
        HCIADD[27]) );
    zao22b U134 ( .A(QHCIADD1[5]), .B(n242), .C(QHCIADD2[5]), .D(n245), .Y(
        HCIADD[5]) );
    zao22b U135 ( .A(QHCIADD1[10]), .B(n242), .C(QHCIADD2[10]), .D(n245), .Y(
        HCIADD[10]) );
    zao22b U136 ( .A(QHCIADD1[25]), .B(n246), .C(QHCIADD2[25]), .D(n266), .Y(
        HCIADD[25]) );
    zivc U137 ( .A(n241), .Y(n269) );
    zivb U138 ( .A(n262), .Y(n247) );
    zivc U139 ( .A(n262), .Y(n252) );
    zivb U140 ( .A(n260), .Y(n248) );
    zao2x4b U141 ( .A(n250), .B(ASYNCLISTADDR[9]), .C(n251), .D(ADI[9]), .E(
        n247), .F(DW1_0[9]), .G(n248), .H(DW2_0[9]), .Y(ASYNCLISTADDR136_9) );
    zao2x4b U142 ( .A(n265), .B(ASYNCLISTADDR[14]), .C(ADI[14]), .D(n251), .E(
        DW1_0[14]), .F(n247), .G(DW2_0[14]), .H(n248), .Y(ASYNCLISTADDR136_14)
         );
    zao2x4b U143 ( .A(n265), .B(ASYNCLISTADDR[20]), .C(ADI[20]), .D(n251), .E(
        DW1_0[20]), .F(n252), .G(DW2_0[20]), .H(n253), .Y(ASYNCLISTADDR136_20)
         );
    zao2x4b U144 ( .A(n265), .B(ASYNCLISTADDR[12]), .C(ADI[12]), .D(n251), .E(
        DW1_0[12]), .F(n252), .G(DW2_0[12]), .H(n253), .Y(ASYNCLISTADDR136_12)
         );
    zao2x4b U145 ( .A(n265), .B(ASYNCLISTADDR[24]), .C(ADI[24]), .D(n251), .E(
        DW1_0[24]), .F(n247), .G(DW2_0[24]), .H(n248), .Y(ASYNCLISTADDR136_24)
         );
    zao2x4b U146 ( .A(n250), .B(ASYNCLISTADDR[5]), .C(ADI[5]), .D(n251), .E(
        DW1_0[5]), .F(n247), .G(DW2_0[5]), .H(n248), .Y(ASYNCLISTADDR136_5) );
    zao2x4b U147 ( .A(n265), .B(ASYNCLISTADDR[26]), .C(ADI[26]), .D(n251), .E(
        DW1_0[26]), .F(n247), .G(DW2_0[26]), .H(n248), .Y(ASYNCLISTADDR136_26)
         );
    zao2x4b U148 ( .A(n265), .B(ASYNCLISTADDR[30]), .C(ADI[30]), .D(n251), .E(
        DW1_0[30]), .F(n252), .G(DW2_0[30]), .H(n253), .Y(ASYNCLISTADDR136_30)
         );
    zao2x4b U149 ( .A(n265), .B(ASYNCLISTADDR[22]), .C(ADI[22]), .D(n251), .E(
        DW1_0[22]), .F(n252), .G(DW2_0[22]), .H(n253), .Y(ASYNCLISTADDR136_22)
         );
    zao2x4b U150 ( .A(n265), .B(ASYNCLISTADDR[10]), .C(ADI[10]), .D(n251), .E(
        DW1_0[10]), .F(n247), .G(DW2_0[10]), .H(n248), .Y(ASYNCLISTADDR136_10)
         );
    zao2x4b U151 ( .A(n250), .B(ASYNCLISTADDR[7]), .C(ADI[7]), .D(n251), .E(
        DW1_0[7]), .F(n247), .G(DW2_0[7]), .H(n248), .Y(ASYNCLISTADDR136_7) );
    zao2x4b U152 ( .A(n265), .B(ASYNCLISTADDR[18]), .C(ADI[18]), .D(n251), .E(
        DW1_0[18]), .F(n252), .G(DW2_0[18]), .H(n253), .Y(ASYNCLISTADDR136_18)
         );
    zao2x4b U153 ( .A(n265), .B(ASYNCLISTADDR[28]), .C(ADI[28]), .D(n251), .E(
        DW1_0[28]), .F(n247), .G(DW2_0[28]), .H(n248), .Y(ASYNCLISTADDR136_28)
         );
    zao2x4b U154 ( .A(n265), .B(ASYNCLISTADDR[16]), .C(ADI[16]), .D(n251), .E(
        DW1_0[16]), .F(n252), .G(DW2_0[16]), .H(n253), .Y(ASYNCLISTADDR136_16)
         );
    zao2x4b U155 ( .A(n250), .B(ASYNCLISTADDR[17]), .C(ADI[17]), .D(
        ASYNCADDR_WE), .E(DW1_0[17]), .F(n252), .G(DW2_0[17]), .H(n253), .Y(
        ASYNCLISTADDR136_17) );
    zao2x4b U156 ( .A(n250), .B(ASYNCLISTADDR[25]), .C(ADI[25]), .D(
        ASYNCADDR_WE), .E(DW1_0[25]), .F(n252), .G(DW2_0[25]), .H(n253), .Y(
        ASYNCLISTADDR136_25) );
    zao2x4b U157 ( .A(n250), .B(ASYNCLISTADDR[19]), .C(ADI[19]), .D(
        ASYNCADDR_WE), .E(DW1_0[19]), .F(n252), .G(DW2_0[19]), .H(n253), .Y(
        ASYNCLISTADDR136_19) );
    zao2x4b U158 ( .A(n265), .B(ASYNCLISTADDR[6]), .C(ADI[6]), .D(ASYNCADDR_WE
        ), .E(DW1_0[6]), .F(n252), .G(DW2_0[6]), .H(n253), .Y(
        ASYNCLISTADDR136_6) );
    zao2x4b U159 ( .A(n250), .B(ASYNCLISTADDR[31]), .C(ADI[31]), .D(
        ASYNCADDR_WE), .E(DW1_0[31]), .F(n252), .G(DW2_0[31]), .H(n253), .Y(
        ASYNCLISTADDR136_31) );
    zao2x4b U160 ( .A(n250), .B(ASYNCLISTADDR[11]), .C(ADI[11]), .D(
        ASYNCADDR_WE), .E(DW1_0[11]), .F(n252), .G(DW2_0[11]), .H(n253), .Y(
        ASYNCLISTADDR136_11) );
    zao2x4b U161 ( .A(n250), .B(ASYNCLISTADDR[29]), .C(ADI[29]), .D(
        ASYNCADDR_WE), .E(DW1_0[29]), .F(n252), .G(DW2_0[29]), .H(n253), .Y(
        ASYNCLISTADDR136_29) );
    zao2x4b U162 ( .A(n250), .B(ASYNCLISTADDR[23]), .C(ADI[23]), .D(
        ASYNCADDR_WE), .E(DW1_0[23]), .F(n252), .G(DW2_0[23]), .H(n253), .Y(
        ASYNCLISTADDR136_23) );
    zao2x4b U163 ( .A(n250), .B(ASYNCLISTADDR[27]), .C(ADI[27]), .D(
        ASYNCADDR_WE), .E(DW1_0[27]), .F(n252), .G(DW2_0[27]), .H(n253), .Y(
        ASYNCLISTADDR136_27) );
    zao2x4b U164 ( .A(n250), .B(ASYNCLISTADDR[13]), .C(ADI[13]), .D(
        ASYNCADDR_WE), .E(DW1_0[13]), .F(n252), .G(DW2_0[13]), .H(n253), .Y(
        ASYNCLISTADDR136_13) );
    zao2x4b U165 ( .A(n250), .B(ASYNCLISTADDR[21]), .C(ADI[21]), .D(
        ASYNCADDR_WE), .E(DW1_0[21]), .F(n252), .G(DW2_0[21]), .H(n253), .Y(
        ASYNCLISTADDR136_21) );
    zao2x4b U166 ( .A(n265), .B(ASYNCLISTADDR[8]), .C(ADI[8]), .D(ASYNCADDR_WE
        ), .E(DW1_0[8]), .F(n252), .G(DW2_0[8]), .H(n253), .Y(
        ASYNCLISTADDR136_8) );
    zao2x4b U167 ( .A(n250), .B(ASYNCLISTADDR[15]), .C(ADI[15]), .D(
        ASYNCADDR_WE), .E(DW1_0[15]), .F(n252), .G(DW2_0[15]), .H(n253), .Y(
        ASYNCLISTADDR136_15) );
    zivc U168 ( .A(n260), .Y(n253) );
    zxo2b U169 ( .A(add_50_carry_29), .B(HCIADR_p_29), .Y(HCIADR[31]) );
    zan2b U170 ( .A(HCIADR_p_28), .B(add_50_carry_28), .Y(add_50_carry_29) );
    zxo2b U171 ( .A(HCIADR_p_28), .B(add_50_carry_28), .Y(HCIADR[30]) );
    zan2b U172 ( .A(HCIADR_p_27), .B(add_50_carry_27), .Y(add_50_carry_28) );
    zxo2b U173 ( .A(HCIADR_p_27), .B(add_50_carry_27), .Y(HCIADR[29]) );
    zan2b U174 ( .A(HCIADR_p_26), .B(add_50_carry_26), .Y(add_50_carry_27) );
    zxo2b U175 ( .A(HCIADR_p_26), .B(add_50_carry_26), .Y(HCIADR[28]) );
    zan2b U176 ( .A(HCIADR_p_25), .B(add_50_carry_25), .Y(add_50_carry_26) );
    zxo2b U177 ( .A(HCIADR_p_25), .B(add_50_carry_25), .Y(HCIADR[27]) );
    zan2b U178 ( .A(HCIADR_p_24), .B(add_50_carry_24), .Y(add_50_carry_25) );
    zxo2b U179 ( .A(HCIADR_p_24), .B(add_50_carry_24), .Y(HCIADR[26]) );
    zan2b U180 ( .A(HCIADR_p_23), .B(add_50_carry_23), .Y(add_50_carry_24) );
    zxo2b U181 ( .A(HCIADR_p_23), .B(add_50_carry_23), .Y(HCIADR[25]) );
    zan2b U182 ( .A(HCIADR_p_22), .B(add_50_carry_22), .Y(add_50_carry_23) );
    zxo2b U183 ( .A(HCIADR_p_22), .B(add_50_carry_22), .Y(HCIADR[24]) );
    zan2b U184 ( .A(HCIADR_p_21), .B(add_50_carry_21), .Y(add_50_carry_22) );
    zxo2b U185 ( .A(HCIADR_p_21), .B(add_50_carry_21), .Y(HCIADR[23]) );
    zan2b U186 ( .A(HCIADR_p_20), .B(add_50_carry_20), .Y(add_50_carry_21) );
    zxo2b U187 ( .A(HCIADR_p_20), .B(add_50_carry_20), .Y(HCIADR[22]) );
    zan2b U188 ( .A(HCIADR_p_19), .B(add_50_carry_19), .Y(add_50_carry_20) );
    zxo2b U189 ( .A(HCIADR_p_19), .B(add_50_carry_19), .Y(HCIADR[21]) );
    zan2b U190 ( .A(HCIADR_p_18), .B(add_50_carry_18), .Y(add_50_carry_19) );
    zxo2b U191 ( .A(HCIADR_p_18), .B(add_50_carry_18), .Y(HCIADR[20]) );
    zan2b U192 ( .A(HCIADR_p_17), .B(add_50_carry_17), .Y(add_50_carry_18) );
    zxo2b U193 ( .A(HCIADR_p_17), .B(add_50_carry_17), .Y(HCIADR[19]) );
    zan2b U194 ( .A(HCIADR_p_16), .B(add_50_carry_16), .Y(add_50_carry_17) );
    zxo2b U195 ( .A(HCIADR_p_16), .B(add_50_carry_16), .Y(HCIADR[18]) );
    zan2b U196 ( .A(HCIADR_p_15), .B(add_50_carry_15), .Y(add_50_carry_16) );
    zxo2b U197 ( .A(HCIADR_p_15), .B(add_50_carry_15), .Y(HCIADR[17]) );
    zan2b U198 ( .A(HCIADR_p_14), .B(add_50_carry_14), .Y(add_50_carry_15) );
    zxo2b U199 ( .A(HCIADR_p_14), .B(add_50_carry_14), .Y(HCIADR[16]) );
    zan2b U200 ( .A(HCIADR_p_13), .B(add_50_carry_13), .Y(add_50_carry_14) );
    zxo2b U201 ( .A(HCIADR_p_13), .B(add_50_carry_13), .Y(HCIADR[15]) );
    zan2b U202 ( .A(HCIADR_p_12), .B(add_50_carry_12), .Y(add_50_carry_13) );
    zxo2b U203 ( .A(HCIADR_p_12), .B(add_50_carry_12), .Y(HCIADR[14]) );
    zan2b U204 ( .A(HCIADR_p_11), .B(add_50_carry_11), .Y(add_50_carry_12) );
    zxo2b U205 ( .A(HCIADR_p_11), .B(add_50_carry_11), .Y(HCIADR[13]) );
    zan2b U206 ( .A(HCIADR_p_10), .B(add_50_carry_10), .Y(add_50_carry_11) );
    zxo2b U207 ( .A(HCIADR_p_10), .B(add_50_carry_10), .Y(HCIADR[12]) );
    zan2b U208 ( .A(HCIADR_p_9), .B(add_50_carry_9), .Y(add_50_carry_10) );
    zxo2b U209 ( .A(HCIADR_p_9), .B(add_50_carry_9), .Y(HCIADR[11]) );
    zan2b U210 ( .A(HCIADR_p_8), .B(add_50_carry_8), .Y(add_50_carry_9) );
    zxo2b U211 ( .A(HCIADR_p_8), .B(add_50_carry_8), .Y(HCIADR[10]) );
    zan2b U212 ( .A(HCIADR_p_7), .B(add_50_carry_7), .Y(add_50_carry_8) );
    zxo2b U213 ( .A(HCIADR_p_7), .B(add_50_carry_7), .Y(HCIADR[9]) );
    zan2b U214 ( .A(HCIADR_p_6), .B(add_50_carry_6), .Y(add_50_carry_7) );
    zxo2b U215 ( .A(HCIADR_p_6), .B(add_50_carry_6), .Y(HCIADR[8]) );
    zan2b U216 ( .A(HCIADR_p_5), .B(add_50_carry_5), .Y(add_50_carry_6) );
    zxo2b U217 ( .A(HCIADR_p_5), .B(add_50_carry_5), .Y(HCIADR[7]) );
    zan2b U218 ( .A(HCIADR_p_4), .B(add_50_carry_4), .Y(add_50_carry_5) );
    zxo2b U219 ( .A(HCIADR_p_4), .B(add_50_carry_4), .Y(HCIADR[6]) );
    zan2b U220 ( .A(DWCNT[0]), .B(HCIADR_p_0), .Y(add_50_carry_1) );
    zxo2b U221 ( .A(DWCNT[0]), .B(HCIADR_p_0), .Y(HCIADR[2]) );
    zfa1b add_50_U1_3 ( .A(HCIADR_p_3), .B(DWCNT[3]), .CI(add_50_carry_3), 
        .CO(add_50_carry_4), .S(HCIADR[5]) );
    zfa1b add_50_U1_2 ( .A(HCIADR_p_2), .B(DWCNT[2]), .CI(add_50_carry_2), 
        .CO(add_50_carry_3), .S(HCIADR[4]) );
    zfa1b add_50_U1_1 ( .A(HCIADR_p_1), .B(DWCNT[1]), .CI(add_50_carry_1), 
        .CO(add_50_carry_2), .S(HCIADR[3]) );
    zao222b U222 ( .A(QHCIADR1[2]), .B(n246), .C(QHCIADR2[2]), .D(n245), .E(
        ASYNCLISTADDR[2]), .F(n270), .Y(HCIADR_p_0) );
    zao222b U223 ( .A(QHCIADR1[3]), .B(n242), .C(QHCIADR2[3]), .D(n266), .E(
        ASYNCLISTADDR[3]), .F(n249), .Y(HCIADR_p_1) );
    zao222b U224 ( .A(QHCIADR1[4]), .B(n242), .C(QHCIADR2[4]), .D(n266), .E(
        ASYNCLISTADDR[4]), .F(n270), .Y(HCIADR_p_2) );
    zao222b U225 ( .A(QHCIADR1[5]), .B(n269), .C(QHCIADR2[5]), .D(n267), .E(
        ASYNCLISTADDR[5]), .F(n249), .Y(HCIADR_p_3) );
    zao222b U226 ( .A(QHCIADR1[6]), .B(n269), .C(QHCIADR2[6]), .D(n267), .E(
        ASYNCLISTADDR[6]), .F(n270), .Y(HCIADR_p_4) );
    zao222b U227 ( .A(QHCIADR1[7]), .B(n242), .C(QHCIADR2[7]), .D(n267), .E(
        ASYNCLISTADDR[7]), .F(n249), .Y(HCIADR_p_5) );
    zao222b U228 ( .A(QHCIADR1[8]), .B(n269), .C(QHCIADR2[8]), .D(n244), .E(
        ASYNCLISTADDR[8]), .F(n270), .Y(HCIADR_p_6) );
    zao222b U229 ( .A(QHCIADR1[9]), .B(n242), .C(QHCIADR2[9]), .D(n267), .E(
        ASYNCLISTADDR[9]), .F(n249), .Y(HCIADR_p_7) );
    zao222b U230 ( .A(QHCIADR1[10]), .B(n269), .C(QHCIADR2[10]), .D(n267), .E(
        ASYNCLISTADDR[10]), .F(n270), .Y(HCIADR_p_8) );
    zao222b U231 ( .A(QHCIADR1[11]), .B(n269), .C(QHCIADR2[11]), .D(n244), .E(
        n249), .F(ASYNCLISTADDR[11]), .Y(HCIADR_p_9) );
    zao222b U232 ( .A(QHCIADR1[12]), .B(n246), .C(QHCIADR2[12]), .D(n267), .E(
        ASYNCLISTADDR[12]), .F(n249), .Y(HCIADR_p_10) );
    zao222b U233 ( .A(QHCIADR1[13]), .B(n269), .C(QHCIADR2[13]), .D(n245), .E(
        ASYNCLISTADDR[13]), .F(n270), .Y(HCIADR_p_11) );
    zao222b U234 ( .A(QHCIADR1[14]), .B(n242), .C(QHCIADR2[14]), .D(n267), .E(
        ASYNCLISTADDR[14]), .F(n249), .Y(HCIADR_p_12) );
    zao222b U235 ( .A(QHCIADR1[15]), .B(n242), .C(QHCIADR2[15]), .D(n267), .E(
        ASYNCLISTADDR[15]), .F(n270), .Y(HCIADR_p_13) );
    zao222b U236 ( .A(QHCIADR1[16]), .B(n269), .C(QHCIADR2[16]), .D(n245), .E(
        ASYNCLISTADDR[16]), .F(n249), .Y(HCIADR_p_14) );
    zao222b U237 ( .A(QHCIADR1[17]), .B(n242), .C(QHCIADR2[17]), .D(n267), .E(
        ASYNCLISTADDR[17]), .F(n270), .Y(HCIADR_p_15) );
    zao222b U238 ( .A(QHCIADR1[18]), .B(n246), .C(QHCIADR2[18]), .D(n267), .E(
        ASYNCLISTADDR[18]), .F(n249), .Y(HCIADR_p_16) );
    zao222b U239 ( .A(QHCIADR1[19]), .B(n269), .C(QHCIADR2[19]), .D(n267), .E(
        ASYNCLISTADDR[19]), .F(n270), .Y(HCIADR_p_17) );
    zao222b U240 ( .A(QHCIADR1[20]), .B(n269), .C(QHCIADR2[20]), .D(n267), .E(
        ASYNCLISTADDR[20]), .F(n249), .Y(HCIADR_p_18) );
    zao222b U241 ( .A(QHCIADR1[21]), .B(n242), .C(QHCIADR2[21]), .D(n266), .E(
        ASYNCLISTADDR[21]), .F(n270), .Y(HCIADR_p_19) );
    zao222b U242 ( .A(QHCIADR1[22]), .B(n242), .C(QHCIADR2[22]), .D(n267), .E(
        ASYNCLISTADDR[22]), .F(n249), .Y(HCIADR_p_20) );
    zao222b U243 ( .A(QHCIADR1[23]), .B(n246), .C(QHCIADR2[23]), .D(n267), .E(
        ASYNCLISTADDR[23]), .F(n270), .Y(HCIADR_p_21) );
    zao222b U244 ( .A(QHCIADR1[24]), .B(n246), .C(QHCIADR2[24]), .D(n244), .E(
        ASYNCLISTADDR[24]), .F(n249), .Y(HCIADR_p_22) );
    zao222b U245 ( .A(QHCIADR1[25]), .B(n246), .C(QHCIADR2[25]), .D(n245), .E(
        ASYNCLISTADDR[25]), .F(n270), .Y(HCIADR_p_23) );
    zao222b U246 ( .A(QHCIADR1[26]), .B(n246), .C(QHCIADR2[26]), .D(n244), .E(
        ASYNCLISTADDR[26]), .F(n249), .Y(HCIADR_p_24) );
    zao222b U247 ( .A(QHCIADR1[27]), .B(n269), .C(QHCIADR2[27]), .D(n266), .E(
        ASYNCLISTADDR[27]), .F(n270), .Y(HCIADR_p_25) );
    zao222b U248 ( .A(QHCIADR1[28]), .B(n246), .C(QHCIADR2[28]), .D(n244), .E(
        ASYNCLISTADDR[28]), .F(n249), .Y(HCIADR_p_26) );
    zao222b U249 ( .A(QHCIADR1[29]), .B(n246), .C(QHCIADR2[29]), .D(n267), .E(
        ASYNCLISTADDR[29]), .F(n270), .Y(HCIADR_p_27) );
    zao222b U250 ( .A(QHCIADR1[30]), .B(n246), .C(QHCIADR2[30]), .D(n266), .E(
        ASYNCLISTADDR[30]), .F(n249), .Y(HCIADR_p_28) );
    zao222b U251 ( .A(QHCIADR1[31]), .B(n242), .C(QHCIADR2[31]), .D(n245), .E(
        ASYNCLISTADDR[31]), .F(n270), .Y(HCIADR_p_29) );
    zoa21d U252 ( .A(ASYNC_ACT), .B(ASYNC_EN), .C(RUN), .Y(n254) );
    zoa21d U253 ( .A(ASYNC_EMPTY2), .B(n256), .C(n257), .Y(n255) );
    zor5b U254 ( .A(n261), .B(ASYNC_EMPTY2), .C(n256), .D(n259), .E(n251), .Y(
        n260) );
    zind2d U255 ( .A(ASYNC_EMPTY1), .B(PARSEQHEND1), .Y(n257) );
    zor3b U256 ( .A(n257), .B(n259), .C(ASYNCADDR_WE), .Y(n262) );
    zind2d U257 ( .A(n254), .B(WR_ASYNCADDR), .Y(n263) );
endmodule


module EHCIFLOW ( PCIDMA_SEL, USBDMA_SEL, LIST_SEL, ASYNC_EXE1, ASYNC_EXE2, 
    PER_EXE1, PER_EXE2, CREQ1, CREQ2, CREQ3, CREQ4, ASYNC_EN, PERIOD_EN, 
    SOFGEN, PRESOF, EOF1, EOF2, FRNUM, PRESOF_EVAL, HCI_PRESOF, PERIOD_PRESOF, 
    TXSOF, EHCI_MAC_EOT, PER_CMDSTART_REQ1, PER_CMDSTART_REQ2, 
    ASYNC_CMDSTART_REQ1, ASYNC_CMDSTART_REQ2, EN_DBG_PORT, DBG_CMDSTART_REQ, 
    DBG_CMDSTART, DBG_ACT, ASYNC_ACT, DBG_LIST, PERIOD_END, PER_CMDSTART1, 
    PER_CMDSTART2, ASYNC_CMDSTART1, ASYNC_CMDSTART2, TCMDSTART, TEST_PACKET, 
    SLAVEMODE, SLCMDSTART, CMDSTART, RUN, SWDBG, EHCIFLOW_IDLE, CLK60M, PCICLK, 
    TRST_ );
output [3:0] PCIDMA_SEL;
output [4:0] USBDMA_SEL;
input  [13:0] FRNUM;
input  ASYNC_EXE1, ASYNC_EXE2, PER_EXE1, PER_EXE2, CREQ1, CREQ2, CREQ3, CREQ4, 
    ASYNC_EN, PERIOD_EN, SOFGEN, PRESOF, EOF1, EOF2, TXSOF, EHCI_MAC_EOT, 
    PER_CMDSTART_REQ1, PER_CMDSTART_REQ2, ASYNC_CMDSTART_REQ1, 
    ASYNC_CMDSTART_REQ2, EN_DBG_PORT, DBG_CMDSTART_REQ, DBG_ACT, ASYNC_ACT, 
    PERIOD_END, TCMDSTART, TEST_PACKET, SLAVEMODE, SLCMDSTART, RUN, SWDBG, 
    CLK60M, PCICLK, TRST_;
output LIST_SEL, PRESOF_EVAL, HCI_PRESOF, PERIOD_PRESOF, DBG_CMDSTART, 
    DBG_LIST, PER_CMDSTART1, PER_CMDSTART2, ASYNC_CMDSTART1, ASYNC_CMDSTART2, 
    CMDSTART, EHCIFLOW_IDLE;
    wire EHCISM_1, CMDSTART_REQ, SPAREO6, USBDMA_SEL642_4, CMDSTART_REQ_PRE, 
        PERIOD_RUN_FIRST975, PERIOD_RUN, SPAREO0_, SPAREO8, PER_TOKEN, 
        W4SOFGEN, CMDREQ_T, PCIDMA_SEL452_2, USBDMA_SEL642_3, EHCISMNXT_1, 
        SPAREO1, CMDSTART_NORM, SPAREO9, EHCISMNXT_0, SPAREO0, USBDMA_SEL642_2, 
        PCIDMA_SEL452_3, EHCISM_0, SPAREO7, val616_1, EOFSOF_P, val540_1, 
        TXSOF_T, CMDSTART_NORM1238, EHCISM_2, SPAREO5, EOFSOF, CMDREQ1164, 
        ASYNC_TOKEN, PCIDMA_SEL452_1, USBDMA_SEL642_0, SPAREO2, EHCISMNXT_2, 
        W4SOFGEN810, SPAREO3, SPAREO1_, EHCISMNXT_3, USBDMA_SEL642_1, 
        PCIDMA_SEL452_0, EHCISM_3, SPAREO4, EOF1_PCLK, n1349, n1350, n1351, 
        n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, 
        n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, 
        n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, 
        n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
        n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
        n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
        n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, 
        n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, 
        n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, 
        n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, 
        n1452, n1453, n1454, n1455, n1456;
    znd3b SPARE519 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE510 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE517 ( .A(SPAREO4), .Y(SPAREO5) );
    znr3b SPARE516 ( .A(SPAREO2), .B(CMDSTART_REQ_PRE), .C(SPAREO0_), .Y(
        SPAREO4) );
    zivb SPARE518 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE511 ( .CK(CLK60M), .D(SPAREO7), .R(TRST_), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zaoi211b SPARE513 ( .A(SPAREO4), .B(EOFSOF_P), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zoai21b SPARE514 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zoai21b SPARE515 ( .A(SPAREO1), .B(DBG_LIST), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE512 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zor2b U340 ( .A(EOF2), .B(SOFGEN), .Y(EOFSOF_P) );
    zmux21lb U341 ( .A(n1358), .B(n1357), .S(n1401), .Y(n1400) );
    zmux21lb U342 ( .A(n1403), .B(n1402), .S(LIST_SEL), .Y(n1401) );
    zor2b U343 ( .A(n1425), .B(n1426), .Y(n1424) );
    zmux21lb U344 ( .A(n1419), .B(n1421), .S(n1359), .Y(n1425) );
    zmux21lb U345 ( .A(n1416), .B(n1418), .S(n1359), .Y(n1426) );
    zor2b U346 ( .A(n1357), .B(n1358), .Y(n1423) );
    zivb U347 ( .A(n1423), .Y(n1422) );
    zmux21lb U348 ( .A(n1444), .B(n1443), .S(LIST_SEL), .Y(n1445) );
    zan2b U349 ( .A(n1349), .B(n1437), .Y(n1444) );
    zan2b U350 ( .A(n1350), .B(n1424), .Y(n1443) );
    zmux21lb U351 ( .A(n1442), .B(n1441), .S(LIST_SEL), .Y(n1446) );
    zan2b U352 ( .A(n1349), .B(n1400), .Y(n1442) );
    zan2b U353 ( .A(n1350), .B(n1435), .Y(n1441) );
    znr4b U354 ( .A(FRNUM[0]), .B(FRNUM[1]), .C(FRNUM[2]), .D(n1398), .Y(n1397
        ) );
    zmux21lb U355 ( .A(n1434), .B(n1433), .S(LIST_SEL), .Y(n1440) );
    zan2b U356 ( .A(n1350), .B(n1435), .Y(n1434) );
    zivb U357 ( .A(n1424), .Y(n1435) );
    zan2b U358 ( .A(n1349), .B(n1400), .Y(n1433) );
    zmux21lb U359 ( .A(n1438), .B(n1436), .S(LIST_SEL), .Y(n1439) );
    zan2b U360 ( .A(n1350), .B(n1424), .Y(n1438) );
    zan2b U361 ( .A(n1349), .B(n1437), .Y(n1436) );
    zivb U362 ( .A(n1400), .Y(n1437) );
    zor2b U363 ( .A(EHCISM_3), .B(EHCISM_0), .Y(n1404) );
    zao32b U364 ( .A(n1352), .B(n1388), .C(n1431), .D(n1351), .E(n1409), .Y(
        n1399) );
    zivb U365 ( .A(DBG_ACT), .Y(n1409) );
    zor2b U366 ( .A(EHCISM_2), .B(EHCISM_1), .Y(n1407) );
    zan2b U367 ( .A(SLAVEMODE), .B(SLCMDSTART), .Y(n1447) );
    zan2b U368 ( .A(USBDMA_SEL[0]), .B(PER_CMDSTART_REQ1), .Y(n1360) );
    zor2b U369 ( .A(TXSOF), .B(TXSOF_T), .Y(n1366) );
    zivb U370 ( .A(n1452), .Y(n1454) );
    zivb U371 ( .A(PRESOF), .Y(n1369) );
    zan2b U372 ( .A(PCIDMA_SEL[1]), .B(n1372), .Y(n1375) );
    zmux21lb U373 ( .A(n1445), .B(n1446), .S(PER_TOKEN), .Y(n1376) );
    zoai2x4b U374 ( .A(n1421), .B(n1387), .C(n1419), .D(n1420), .E(n1418), .F(
        n1371), .G(n1416), .H(n1417), .Y(n1372) );
    zivb U375 ( .A(CREQ3), .Y(n1421) );
    zivb U376 ( .A(CREQ4), .Y(n1419) );
    zivb U377 ( .A(CREQ1), .Y(n1418) );
    zivb U378 ( .A(CREQ2), .Y(n1416) );
    zivb U379 ( .A(n1428), .Y(n1427) );
    zmux21lb U380 ( .A(n1446), .B(n1445), .S(PER_TOKEN), .Y(n1374) );
    zan2b U381 ( .A(n1384), .B(n1385), .Y(n1383) );
    zan2b U382 ( .A(ASYNC_EXE1), .B(n1353), .Y(USBDMA_SEL642_2) );
    zor2b U383 ( .A(EHCISMNXT_0), .B(n1386), .Y(n1370) );
    zmux21lb U384 ( .A(n1440), .B(n1439), .S(ASYNC_TOKEN), .Y(n1378) );
    zivb U385 ( .A(n1372), .Y(n1451) );
    zao32b U386 ( .A(n1388), .B(n1352), .C(n1389), .D(n1351), .E(DBG_ACT), .Y(
        EHCISMNXT_1) );
    zivb U387 ( .A(n1410), .Y(n1388) );
    zivb U388 ( .A(n1431), .Y(n1389) );
    znd2b U389 ( .A(DBG_ACT), .B(EN_DBG_PORT), .Y(n1431) );
    zan2b U390 ( .A(n1356), .B(n1364), .Y(PERIOD_RUN_FIRST975) );
    zan2b U391 ( .A(PCIDMA_SEL[3]), .B(n1372), .Y(n1380) );
    zmux21lb U392 ( .A(n1439), .B(n1440), .S(ASYNC_TOKEN), .Y(n1381) );
    zivb U393 ( .A(TEST_PACKET), .Y(n1377) );
    zan2b U394 ( .A(ASYNC_EXE2), .B(n1353), .Y(USBDMA_SEL642_3) );
    zivb U395 ( .A(n1414), .Y(n1393) );
    zan2b U396 ( .A(n1390), .B(n1452), .Y(n1394) );
    zivb U397 ( .A(n1406), .Y(n1390) );
    zivb U398 ( .A(n1429), .Y(n1395) );
    zivb U399 ( .A(RUN), .Y(n1398) );
    zivb U400 ( .A(n1362), .Y(n1396) );
    zivb U401 ( .A(n1399), .Y(n1412) );
    zor2b U402 ( .A(DBG_LIST), .B(EHCISM_0), .Y(EHCIFLOW_IDLE) );
    zivb U403 ( .A(EHCIFLOW_IDLE), .Y(n1385) );
    zmux21lb U404 ( .A(n1447), .B(TCMDSTART), .S(TEST_PACKET), .Y(n1382) );
    zan2b U405 ( .A(n1355), .B(USBDMA_SEL[3]), .Y(ASYNC_CMDSTART2) );
    zan2b U406 ( .A(n1355), .B(USBDMA_SEL[2]), .Y(ASYNC_CMDSTART1) );
    zan2b U407 ( .A(n1355), .B(USBDMA_SEL[1]), .Y(PER_CMDSTART2) );
    zan2b U408 ( .A(n1355), .B(USBDMA_SEL[0]), .Y(PER_CMDSTART1) );
    zan2b U409 ( .A(n1355), .B(USBDMA_SEL[4]), .Y(DBG_CMDSTART) );
    zan2b U410 ( .A(CMDSTART_REQ_PRE), .B(n1365), .Y(PRESOF_EVAL) );
    zdffqsb HCI_PRESOF_reg ( .CK(PCICLK), .D(PRESOF), .S(TRST_), .Q(HCI_PRESOF
        ) );
    zivb U411 ( .A(HCI_PRESOF), .Y(n1368) );
    zdffqrb USBDMA_SEL_reg_1 ( .CK(PCICLK), .D(USBDMA_SEL642_1), .R(TRST_), 
        .Q(USBDMA_SEL[1]) );
    zdffqrb CMDSTART_NORM_reg ( .CK(PCICLK), .D(CMDSTART_NORM1238), .R(TRST_), 
        .Q(CMDSTART_NORM) );
    zivb U412 ( .A(CMDSTART_NORM), .Y(n1415) );
    zdffrb EHCISM_reg_2 ( .CK(PCICLK), .D(EHCISMNXT_2), .R(TRST_), .Q(EHCISM_2
        ), .QN(n1405) );
    zdffqrb CMDREQ_reg ( .CK(PCICLK), .D(n1456), .R(TRST_), .Q(CMDSTART_REQ)
         );
    zivb U413 ( .A(CMDSTART_REQ), .Y(n1365) );
    zdffqrb PCIDMA_SEL_reg_1 ( .CK(PCICLK), .D(PCIDMA_SEL452_1), .R(TRST_), 
        .Q(PCIDMA_SEL[1]) );
    zivb U414 ( .A(PCIDMA_SEL[1]), .Y(n1417) );
    zdffqsb PCIDMA_SEL_reg_0 ( .CK(PCICLK), .D(PCIDMA_SEL452_0), .S(TRST_), 
        .Q(PCIDMA_SEL[0]) );
    zivb U415 ( .A(PCIDMA_SEL[0]), .Y(n1371) );
    zdffqrb EHCISM_reg_3 ( .CK(PCICLK), .D(EHCISMNXT_3), .R(TRST_), .Q(
        EHCISM_3) );
    zivb U416 ( .A(EHCISM_3), .Y(n1413) );
    zdffqsb USBDMA_SEL_reg_0 ( .CK(PCICLK), .D(USBDMA_SEL642_0), .S(TRST_), 
        .Q(USBDMA_SEL[0]) );
    zdffqrb ASYNC_TOKEN_reg ( .CK(PCICLK), .D(val616_1), .R(TRST_), .Q(
        ASYNC_TOKEN) );
    zivb U417 ( .A(ASYNC_TOKEN), .Y(n1402) );
    zdffqrb USBDMA_SEL_reg_2 ( .CK(PCICLK), .D(USBDMA_SEL642_2), .R(TRST_), 
        .Q(USBDMA_SEL[2]) );
    zdffqrb EOF1_PCLK_reg ( .CK(PCICLK), .D(EOF1), .R(TRST_), .Q(EOF1_PCLK) );
    zdffqrb EOFSOF_reg ( .CK(PCICLK), .D(SOFGEN), .R(TRST_), .Q(EOFSOF) );
    zdffqrb PERIOD_RUN_reg ( .CK(PCICLK), .D(n1356), .R(TRST_), .Q(PERIOD_RUN)
         );
    zivb U418 ( .A(PERIOD_RUN), .Y(n1364) );
    zdffqrb W4SOFGEN_reg ( .CK(PCICLK), .D(n1455), .R(TRST_), .Q(W4SOFGEN) );
    zivb U419 ( .A(W4SOFGEN), .Y(n1408) );
    zdffqrb EHCISM_reg_1 ( .CK(PCICLK), .D(EHCISMNXT_1), .R(TRST_), .Q(
        EHCISM_1) );
    zivb U420 ( .A(EHCISM_1), .Y(n1411) );
    zdffrb PCIDMA_SEL_reg_2 ( .CK(PCICLK), .D(PCIDMA_SEL452_2), .R(TRST_), .Q(
        PCIDMA_SEL[2]), .QN(n1387) );
    zdffqrb DBG_LIST_reg ( .CK(PCICLK), .D(EHCISMNXT_1), .R(TRST_), .Q(
        DBG_LIST) );
    zdffrb PERIOD_RUN_FIRST_reg ( .CK(PCICLK), .D(PERIOD_RUN_FIRST975), .R(
        TRST_), .QN(n1453) );
    zdffqrb PCIDMA_SEL_reg_3 ( .CK(PCICLK), .D(PCIDMA_SEL452_3), .R(TRST_), 
        .Q(PCIDMA_SEL[3]) );
    zivb U421 ( .A(PCIDMA_SEL[3]), .Y(n1420) );
    zdffqsb EHCISM_reg_0 ( .CK(PCICLK), .D(EHCISMNXT_0), .S(TRST_), .Q(
        EHCISM_0) );
    zivb U422 ( .A(EHCISM_0), .Y(n1386) );
    zdffqrb USBDMA_SEL_reg_4 ( .CK(PCICLK), .D(USBDMA_SEL642_4), .R(TRST_), 
        .Q(USBDMA_SEL[4]) );
    zdffqrb USBDMA_SEL_reg_3 ( .CK(PCICLK), .D(USBDMA_SEL642_3), .R(TRST_), 
        .Q(USBDMA_SEL[3]) );
    zdffqrb PER_TOKEN_reg ( .CK(PCICLK), .D(val540_1), .R(TRST_), .Q(PER_TOKEN
        ) );
    zivb U423 ( .A(PER_TOKEN), .Y(n1403) );
    zdffqrb TXSOF_T_reg ( .CK(PCICLK), .D(TXSOF), .R(TRST_), .Q(TXSOF_T) );
    zdffrb LIST_SEL_reg ( .CK(PCICLK), .D(EHCISMNXT_3), .R(TRST_), .Q(LIST_SEL
        ), .QN(n1384) );
    zdffqrb CMDREQ_T_reg ( .CK(PCICLK), .D(CMDSTART_REQ_PRE), .R(TRST_), .Q(
        CMDREQ_T) );
    znr2b U424 ( .A(n1422), .B(n1372), .Y(n1349) );
    znr3b U425 ( .A(n1427), .B(n1423), .C(n1372), .Y(n1350) );
    znr3b U426 ( .A(EHCISM_2), .B(n1411), .C(n1404), .Y(n1351) );
    znr2b U427 ( .A(EOFSOF), .B(n1408), .Y(n1352) );
    znr3b U428 ( .A(EHCISM_0), .B(n1384), .C(TEST_PACKET), .Y(n1353) );
    zoa211b U429 ( .A(RUN), .B(ASYNC_ACT), .C(n1368), .D(n1430), .Y(n1354) );
    znr3b U430 ( .A(n1415), .B(SLAVEMODE), .C(TEST_PACKET), .Y(n1355) );
    zmux21hb U431 ( .A(PERIOD_RUN), .B(PERIOD_EN), .S(n1397), .Y(n1356) );
    zmux21hb U432 ( .A(CREQ1), .B(CREQ3), .S(LIST_SEL), .Y(n1357) );
    zmux21hb U433 ( .A(CREQ2), .B(CREQ4), .S(LIST_SEL), .Y(n1358) );
    zmux21hb U434 ( .A(ASYNC_TOKEN), .B(PER_TOKEN), .S(LIST_SEL), .Y(n1359) );
    zao211b U435 ( .A(USBDMA_SEL[1]), .B(PER_CMDSTART_REQ2), .C(n1360), .D(
        n1361), .Y(CMDSTART_REQ_PRE) );
    zoai21b U436 ( .A(ASYNC_EN), .B(n1362), .C(n1363), .Y(EHCISMNXT_0) );
    zoa21d U437 ( .A(USBDMA_SEL[0]), .B(USBDMA_SEL[1]), .C(HCI_PRESOF), .Y(
        PERIOD_PRESOF) );
    zao21b U438 ( .A(CMDSTART_NORM), .B(n1366), .C(n1367), .Y(
        CMDSTART_NORM1238) );
    zan4b U439 ( .A(n1368), .B(CMDREQ_T), .C(n1369), .D(CMDSTART_REQ_PRE), .Y(
        CMDREQ1164) );
    zao21b U440 ( .A(W4SOFGEN), .B(n1370), .C(EOFSOF), .Y(W4SOFGEN810) );
    zao21b U441 ( .A(PER_TOKEN), .B(n1371), .C(PCIDMA_SEL[1]), .Y(val540_1) );
    zao211b U442 ( .A(PCIDMA_SEL[0]), .B(n1372), .C(n1373), .D(n1374), .Y(
        PCIDMA_SEL452_0) );
    zoa21d U443 ( .A(n1375), .B(n1376), .C(n1377), .Y(PCIDMA_SEL452_1) );
    zoa21d U444 ( .A(n1378), .B(n1379), .C(n1377), .Y(PCIDMA_SEL452_2) );
    zoa21d U445 ( .A(n1380), .B(n1381), .C(n1377), .Y(PCIDMA_SEL452_3) );
    zind2b U446 ( .A(n1355), .B(n1382), .Y(CMDSTART) );
    zao21b U447 ( .A(n1383), .B(PER_EXE1), .C(TEST_PACKET), .Y(USBDMA_SEL642_0
        ) );
    zan4b U448 ( .A(n1384), .B(n1385), .C(n1377), .D(PER_EXE2), .Y(
        USBDMA_SEL642_1) );
    zan4b U449 ( .A(DBG_LIST), .B(DBG_ACT), .C(n1377), .D(n1386), .Y(
        USBDMA_SEL642_4) );
    zao21b U450 ( .A(ASYNC_TOKEN), .B(n1387), .C(PCIDMA_SEL[3]), .Y(val616_1)
         );
    zao21b U451 ( .A(n1390), .B(n1391), .C(n1392), .Y(EHCISMNXT_2) );
    zao222b U452 ( .A(n1354), .B(n1393), .C(n1394), .D(n1395), .E(ASYNC_EN), 
        .F(n1396), .Y(EHCISMNXT_3) );
    zoa21d U453 ( .A(PERIOD_RUN), .B(n1356), .C(n1399), .Y(n1392) );
    zan4b U454 ( .A(n1386), .B(n1368), .C(CMDSTART_REQ), .D(n1369), .Y(n1367)
         );
    zor3b U455 ( .A(EHCISM_1), .B(n1405), .C(n1404), .Y(n1406) );
    zor3b U456 ( .A(EHCISM_3), .B(n1386), .C(n1407), .Y(n1410) );
    zor3b U457 ( .A(PERIOD_RUN), .B(n1412), .C(n1356), .Y(n1362) );
    zor3b U458 ( .A(EHCISM_0), .B(n1413), .C(n1407), .Y(n1414) );
    zor4b U459 ( .A(CREQ1), .B(CREQ2), .C(CREQ3), .D(CREQ4), .Y(n1428) );
    zor3b U460 ( .A(W4SOFGEN), .B(EOF1_PCLK), .C(n1398), .Y(n1429) );
    zxo2b U461 ( .A(n1407), .B(n1404), .Y(n1432) );
    zoa22b U462 ( .A(n1354), .B(n1414), .C(n1352), .D(n1410), .Y(n1448) );
    zan4b U463 ( .A(n1449), .B(n1432), .C(n1450), .D(n1448), .Y(n1363) );
    zoa22b U464 ( .A(n1405), .B(n1411), .C(n1386), .D(n1413), .Y(n1449) );
    zao222b U465 ( .A(USBDMA_SEL[4]), .B(DBG_CMDSTART_REQ), .C(USBDMA_SEL[3]), 
        .D(ASYNC_CMDSTART_REQ2), .E(USBDMA_SEL[2]), .F(ASYNC_CMDSTART_REQ1), 
        .Y(n1361) );
    zoai22b U466 ( .A(n1451), .B(n1387), .C(n1384), .D(n1428), .Y(n1379) );
    zao21b U467 ( .A(n1427), .B(n1384), .C(TEST_PACKET), .Y(n1373) );
    zao21b U468 ( .A(PERIOD_END), .B(n1453), .C(HCI_PRESOF), .Y(n1452) );
    zoai21b U469 ( .A(EOF1_PCLK), .B(W4SOFGEN), .C(EHCI_MAC_EOT), .Y(n1430) );
    zor4b U470 ( .A(n1395), .B(n1406), .C(SWDBG), .D(n1454), .Y(n1450) );
    zao21b U471 ( .A(SWDBG), .B(n1429), .C(n1454), .Y(n1391) );
    zbfb U472 ( .A(W4SOFGEN810), .Y(n1455) );
    zbfb U473 ( .A(CMDREQ1164), .Y(n1456) );
endmodule


module EHCI_MUX ( GEN_PERR1, GEN_PERR2, GEN_PERR, RUN_C1, RUN_C2, RUN_C, 
    FROZEN1, FROZEN2, FROZEN, TEST_PACKET, SLAVE_ACT, TRST_, ATPG_ENI, 
    BMUCRST_, PER_BUI_GO1, TBUI_GO, SLBUI_GO, SLAVEMODE, BUI_GO1, ITDIOCINT_S1, 
    ITDIOCINT_S2, QHIOCINT_S1, QHIOCINT_S2, QHIOCINT_S3, QHIOCINT_S4, 
    SITDIOCINT_S1, SITDIOCINT_S2, ITDERRINT_S1, ITDERRINT_S2, QHERRINT_S1, 
    QHERRINT_S2, QHERRINT_S3, QHERRINT_S4, SITDERRINT_S1, SITDERRINT_S2, 
    USBINT_S, ERRINT_S, EHCIFLOW_IDLE, ASYNC_ACT, PERIOD_END, EHCI_IDLE );
input  GEN_PERR1, GEN_PERR2, RUN_C1, RUN_C2, FROZEN1, FROZEN2, TEST_PACKET, 
    SLAVE_ACT, TRST_, ATPG_ENI, PER_BUI_GO1, TBUI_GO, SLBUI_GO, SLAVEMODE, 
    ITDIOCINT_S1, ITDIOCINT_S2, QHIOCINT_S1, QHIOCINT_S2, QHIOCINT_S3, 
    QHIOCINT_S4, SITDIOCINT_S1, SITDIOCINT_S2, ITDERRINT_S1, ITDERRINT_S2, 
    QHERRINT_S1, QHERRINT_S2, QHERRINT_S3, QHERRINT_S4, SITDERRINT_S1, 
    SITDERRINT_S2, EHCIFLOW_IDLE, ASYNC_ACT, PERIOD_END;
output GEN_PERR, RUN_C, FROZEN, BMUCRST_, BUI_GO1, USBINT_S, ERRINT_S, 
    EHCI_IDLE;
    wire n269, n270, n271, n272;
    zao21b U24 ( .A(n269), .B(TRST_), .C(ATPG_ENI), .Y(BMUCRST_) );
    zan3b U25 ( .A(PERIOD_END), .B(n270), .C(EHCIFLOW_IDLE), .Y(EHCI_IDLE) );
    zor2b U26 ( .A(RUN_C2), .B(RUN_C1), .Y(RUN_C) );
    zor2b U27 ( .A(GEN_PERR2), .B(GEN_PERR1), .Y(GEN_PERR) );
    zor5b U28 ( .A(ITDERRINT_S1), .B(ITDERRINT_S2), .C(SITDERRINT_S2), .D(
        SITDERRINT_S1), .E(n271), .Y(ERRINT_S) );
    zor5b U29 ( .A(SITDIOCINT_S2), .B(QHIOCINT_S4), .C(ITDIOCINT_S2), .D(
        SITDIOCINT_S1), .E(n272), .Y(USBINT_S) );
    zor2b U30 ( .A(FROZEN2), .B(FROZEN1), .Y(FROZEN) );
    zmux31hb U31 ( .A(SLAVEMODE), .B(TEST_PACKET), .D0(PER_BUI_GO1), .D1(
        SLBUI_GO), .D2(TBUI_GO), .Y(BUI_GO1) );
    zor4b U32 ( .A(QHIOCINT_S3), .B(ITDIOCINT_S1), .C(QHIOCINT_S2), .D(
        QHIOCINT_S1), .Y(n272) );
    zor4b U33 ( .A(QHERRINT_S1), .B(QHERRINT_S3), .C(QHERRINT_S4), .D(
        QHERRINT_S2), .Y(n271) );
    znr2b U34 ( .A(TEST_PACKET), .B(SLAVE_ACT), .Y(n269) );
    zivb U35 ( .A(ASYNC_ACT), .Y(n270) );
endmodule


module PERIODICFLOW ( PERIOD_EN, PCIEND, GEN_PERR, DWNUM, HCI_PRESOF, 
    PHCI_PRESOF, TDSTARTADR, EHCIREQ, RUN, PERIOD_ACT, PARSETDEND1, 
    PARSETDEND2, TD_PARSE_GO1, TD_PARSE_GO2, TDPARSING1, TDPARSING2, 
    PERIOD_END, PCACHE_EN, PHCI_DW0, PHCI_DW1, DW1_0, DW2_0, CACHE_INVALID1, 
    CACHE_INVALID2, EXEITD1, EXEITD2, EXEQH1, EXEQH2, EXESITD1, EXESITD2, 
    ITDIDLE1, ITDIDLE2, QHIDLE1, QHIDLE2, SITDIDLE1, SITDIDLE2, TD_ACT1, 
    TD_ACT2, PER_EXE1, PER_EXE2, TDHCIREQ1, TDHCIREQ2, TDHCIGNT1, TDHCIGNT2, 
    TD_CACHE_EN1, TD_CACHE_EN2, DWOFFSET, PERHCIADR, CACHE_ADDR1, CACHE_ADDR2, 
    CACHE_EN1, CACHE_EN2, LIST_SEL, TDEXE1, TDEXE2, LTINT_PCLK, SWDBG, RUN_C, 
    FROZEN, FRNUM, FRNUM_PER, FLBASE, TDCMDSTART1, TDCMDSTART2, RECOVERYMODE, 
    EHCIFLOW_IDLE, TDIDLE1, TDIDLE2, FRLSTSIZE, PCICLK, TRST_ );
output [3:0] DWNUM;
input  [31:0] DW2_0;
output [26:0] CACHE_ADDR2;
input  [13:0] FRNUM;
input  [1:0] FRLSTSIZE;
output [3:0] DWOFFSET;
output [31:0] TDSTARTADR;
input  [31:0] PHCI_DW0;
input  [31:0] DW1_0;
input  [31:0] PHCI_DW1;
output [31:0] PERHCIADR;
output [26:0] CACHE_ADDR1;
output [13:0] FRNUM_PER;
input  [19:0] FLBASE;
input  PERIOD_EN, PCIEND, GEN_PERR, HCI_PRESOF, RUN, PARSETDEND1, PARSETDEND2, 
    TDPARSING1, TDPARSING2, CACHE_INVALID1, CACHE_INVALID2, ITDIDLE1, ITDIDLE2, 
    QHIDLE1, QHIDLE2, SITDIDLE1, SITDIDLE2, TDHCIREQ1, TDHCIREQ2, LIST_SEL, 
    TDEXE1, TDEXE2, LTINT_PCLK, SWDBG, TDCMDSTART1, TDCMDSTART2, EHCIFLOW_IDLE, 
    PCICLK, TRST_;
output PHCI_PRESOF, EHCIREQ, PERIOD_ACT, TD_PARSE_GO1, TD_PARSE_GO2, 
    PERIOD_END, PCACHE_EN, EXEITD1, EXEITD2, EXEQH1, EXEQH2, EXESITD1, 
    EXESITD2, TD_ACT1, TD_ACT2, PER_EXE1, PER_EXE2, TDHCIGNT1, TDHCIGNT2, 
    TD_CACHE_EN1, TD_CACHE_EN2, CACHE_EN1, CACHE_EN2, RUN_C, FROZEN, 
    RECOVERYMODE, TDIDLE1, TDIDLE2;
    wire PERIOD_RUN_pre, PERIODSM_3, TD_PARSE_GO2_T, CACHE_ADDR21034_8, 
        FRNUM_INC, SAVEPTR_24, SAVEPTR679_28, SAVEPTR_9, CACHE_ADDR21034_23, 
        TDSTARTADR717_27, CACHE_HIT, SPAREO6, SAVEPTR679_2, EXEITD21109, 
        SAVEPTR679_14, FRNUM_PER_PRE574_8, CACHE_ADDR1996_23, SAVEPTR_18, 
        FRNUM_PER_PRE597_3, CACHE_ADDR1996_16, SAVEPTR_0, CACHE_ADDR21034_1, 
        SAVEPTR679_21, TDSTARTADR717_2, FRNUM_PER_PRE574_11, CACHE_ADDR1996_2, 
        DWNUM1434_3, PERIODSMNXT_0, TDSTARTADR717_12, LAT_SAVEPLACE_COND, 
        CACHE_ADDR21034_16, SAVEPTR_11, FRNUM_PER_PRE574_1, SAVEPTR_31, 
        FRNUM_PER_PRE574_6, SAVEPTR_16, PERIOD_RUN, CACHE_ADDR21034_11, 
        SPAREO0_, TDSTARTADR717_15, TDSTARTADR717_5, TDSTARTADR717_29, SPAREO8, 
        CACHE_ADDR1996_5, CACHE_ADDR21034_6, CACHE_ADDR1996_11, 
        FRNUM_PER_PRE597_4, SAVEPTR679_26, SAVEPTR_7, SAVEPTR679_13, 
        CACHE_ADDR1996_24, SAVEPTR679_5, CACHE_ADDR21034_18, TDSTARTADR717_20, 
        CACHE_ADDR21034_24, SPAREO1, SAVEPTR_23, CACHE_ADDR1996_18, 
        CACHE_ADDR21034_7, CACHE_ADDR1996_10, FRNUM_PER_PRE597_5, 
        SAVEPTR679_27, SAVEPTR_6, TDSTARTADR717_4, TDSTARTADR717_28, 
        CACHE_ADDR1996_4, PERIODSMNXT_6, EXE_HALT, CACHE_ADDR21034_10, 
        FRNUM_PER_PRE597_12, TDSTARTADR717_14, FRNUM_PER_PRE_11, SAVEPTR_30, 
        FRNUM_PER_PRE574_7, SAVEPTR_17, SAVEPTR_22, CACHE_ADDR1996_19, 
        PERIODSM_5, PHASENXT_ParseTD, TDSTARTADR717_21, CACHE_ADDR21034_25, 
        SPAREO0, SAVEPTR679_4, CACHE_ADDR21034_19, SAVEPTR679_12, 
        CACHE_ADDR1996_25, SAVEPTR679_15, FRNUM_PER_PRE574_9, 
        CACHE_ADDR1996_22, SAVEPTR_19, SAVEPTR679_3, CACHEHIT1, 
        CACHE_ADDR21034_22, TDSTARTADR717_26, SPAREO7, CACHE_ADDR21034_9, 
        SAVEPTR_25, SAVEPTR679_29, SAVEPTR_8, EXE_HALT_pre, SAVEPTR_10, 
        FRNUM_PER_PRE574_0, TDSTARTADR717_13, CACHE_ADDR21034_17, EXEQH21183, 
        TDSTARTADR717_3, FRNUM_PER_PRE574_10, CACHE_ADDR1996_3, DWNUM1434_2, 
        FRNUM_PER_PRE597_2, CACHE_ADDR1996_17, CACHE_ADDR21034_0, SAVEPTR_1, 
        SAVEPTR679_20, SAVEPTR_27, FRNUM_PER_PRE597_9, CACHE_ADDR1996_8, 
        CACHE_SEL_PRE, PHASE_FetchFSTN, SPAREO5, TDSTARTADR717_24, 
        TDSTARTADR717_8, CACHE_ADDR21034_20, TDSTARTADR717_18, SAVEPTR679_1, 
        CACHE_ADDR1996_20, FETCHTD, SAVEPTR679_30, SAVEPTR679_17, 
        SAVEPTR679_22, SAVEPTR_3, CACHE_ADDR21034_2, FRNUM_PER_PRE597_0, 
        CACHE_ADDR1996_15, DWNUM1434_0, FRNUM_PER_PRE574_12, CACHE_ADDR1996_1, 
        TDSTARTADR717_1, CACHE_ADDR21034_15, EXESITD11220, TDSTARTADR717_11, 
        SAVEPTR679_8, FRNUM_PER_PRE574_2, SAVEPTR_12, SAVEPTR_15, 
        FRNUM_PER_PRE574_5, SAVEPTR679_19, FRNUM_PER_PRE597_10, 
        TDSTARTADR717_16, TDSTARTADR717_31, CACHE_ADDR21034_12, 
        CACHE_ADDR1996_6, TDSTARTADR717_6, RECOVERYMODE642, SAVEPTR_4, 
        SAVEPTR679_25, CACHE_ADDR1996_12, FRNUM_PER_PRE597_7, SAVEPTR_29, 
        CACHE_ADDR21034_5, TRANEXED1556, SAVEPTR679_10, EXEITD11072, 
        SAVEPTR679_6, FETCHTDNXT, SPAREO2, TDSTARTADR717_23, SAVEPTR_20, 
        CACHE_SEL, SAVEPTR_5, SAVEPTR679_24, CACHE_ADDR1996_13, 
        FRNUM_PER_PRE597_6, SAVEPTR_28, CACHE_ADDR21034_4, CACHE_ADDR1996_7, 
        TDSTARTADR717_7, PHASENXT_FetchTD, FRNUM_PER_PRE597_11, 
        TDSTARTADR717_17, PERIODSM_6, TDSTARTADR717_30, CACHE_ADDR21034_13, 
        PERIODSMNXT_5, SAVEPTR_14, TD_PARSE_GO1_T, FRNUM_PER_PRE574_4, 
        FRNUM_PER_PRE_12, PHASE_ParseTD, SAVEPTR679_18, EXEQH11146, 
        PHASENXT_FetchPList, SAVEPTR_21, SPAREO3, SPAREO1_, CACHE_ADDR21034_26, 
        TDSTARTADR717_22, SAVEPTR679_7, CACHE_ADDR1996_26, SAVEPTR679_11, 
        CACHE_ADDR1996_21, TD_ACT_SEL827, SAVEPTR679_31, SAVEPTR679_16, 
        TDSTARTADR717_19, CACHEHIT2, SAVEPTR679_0, CACHE_ADDR1996_9, 
        PERIODSM_1, SPAREO4, TDSTARTADR717_25, TDSTARTADR717_9, 
        CACHE_ADDR21034_21, EXESITD21257, FRNUM_PER_PRE597_8, SAVEPTR_26, 
        FRNUM_PER_PRE574_3, SAVEPTR_13, FRNUM_INC506, CACHE_ADDR21034_14, 
        TDSTARTADR717_10, SAVEPTR679_9, FROZEN1654, DWNUM1434_1, 
        CACHE_ADDR1996_0, TDSTARTADR717_0, SAVEPTR679_23, TRANEXED, SAVEPTR_2, 
        CACHE_ADDR21034_3, FRNUM_PER_PRE597_1, CACHE_ADDR1996_14, n2009, n2010, 
        n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, 
        add_250_carry_8, add_250_carry_12, add_250_carry_6, add_250_carry_7, 
        add_250_carry_9, add_250_carry_2, add_250_carry_11, add_250_carry_5, 
        add_250_carry_10, add_250_carry_4, add_250_carry_3, n2021, n2022, 
        n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
        n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
        n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
        n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
        n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
        n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
        n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
        n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
        n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
        n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
        n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
        n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
        n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
        n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
        n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
        n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
        n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
        n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
        n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
        n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
        n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
        n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
        n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
        n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
        n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
        n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
        n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
        n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
        n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
        n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
        n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
        n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
        n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
        n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
        n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
        n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
        n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
        n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
        n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
        n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
        n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
        n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, 
        n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, 
        n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, 
        n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, 
        n2483;
    assign DWOFFSET[3] = 1'b0;
    assign DWOFFSET[2] = 1'b0;
    assign DWOFFSET[1] = 1'b0;
    assign DWOFFSET[0] = 1'b0;
    assign PERHCIADR[1] = 1'b0;
    assign PERHCIADR[0] = 1'b0;
    assign FRNUM_PER[13] = 1'b0;
    zdffrb SPARE870 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE879 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb SPARE877 ( .A(SPAREO4), .Y(SPAREO5) );
    znr3b SPARE876 ( .A(SPAREO2), .B(FETCHTD), .C(SPAREO0_), .Y(SPAREO4) );
    zdffrb SPARE871 ( .CK(PCICLK), .D(SPAREO7), .R(TRST_), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE878 ( .A(SPAREO5), .Y(SPAREO6) );
    zaoi211b SPARE873 ( .A(SPAREO4), .B(CACHEHIT2), .C(SPAREO6), .D(
        PERIOD_RUN_pre), .Y(SPAREO8) );
    zoai21b SPARE874 ( .A(SPAREO0), .B(SPAREO8), .C(LAT_SAVEPLACE_COND) );
    zoai21b SPARE875 ( .A(SPAREO1), .B(EXE_HALT_pre), .C(CACHE_HIT), .Y(
        SPAREO3) );
    zaoi211b SPARE872 ( .A(SPAREO0), .B(CACHEHIT1), .C(SPAREO1_), .D(
        FETCHTDNXT), .Y(SPAREO2) );
    zxo2b U745 ( .A(n2209), .B(TDSTARTADR[9]), .Y(n2431) );
    zxo2b U746 ( .A(n2208), .B(TDSTARTADR[29]), .Y(n2432) );
    zxo2b U747 ( .A(n2207), .B(TDSTARTADR[30]), .Y(n2433) );
    zxo2b U748 ( .A(n2212), .B(TDSTARTADR[22]), .Y(n2444) );
    zxo2b U749 ( .A(n2210), .B(TDSTARTADR[14]), .Y(n2443) );
    zxo2b U750 ( .A(n2211), .B(TDSTARTADR[20]), .Y(n2442) );
    zxo2b U751 ( .A(n2216), .B(TDSTARTADR[26]), .Y(n2435) );
    zxo2b U752 ( .A(n2215), .B(TDSTARTADR[8]), .Y(n2436) );
    zxo2b U753 ( .A(n2214), .B(TDSTARTADR[28]), .Y(n2437) );
    zxo2b U754 ( .A(n2213), .B(TDSTARTADR[13]), .Y(n2438) );
    zxo2b U755 ( .A(n2219), .B(TDSTARTADR[25]), .Y(n2441) );
    zxo2b U756 ( .A(n2217), .B(TDSTARTADR[5]), .Y(n2440) );
    zxo2b U757 ( .A(n2218), .B(TDSTARTADR[6]), .Y(n2439) );
    zxo2b U758 ( .A(TDSTARTADR[10]), .B(CACHE_ADDR1[5]), .Y(n2382) );
    zxo2b U759 ( .A(TDSTARTADR[15]), .B(CACHE_ADDR1[10]), .Y(n2383) );
    zxo2b U760 ( .A(TDSTARTADR[27]), .B(CACHE_ADDR1[22]), .Y(n2380) );
    zxo2b U761 ( .A(TDSTARTADR[31]), .B(CACHE_ADDR1[26]), .Y(n2381) );
    zxo2b U762 ( .A(TDSTARTADR[23]), .B(CACHE_ADDR1[18]), .Y(n2386) );
    zxo2b U763 ( .A(TDSTARTADR[24]), .B(CACHE_ADDR1[19]), .Y(n2385) );
    zxo2b U764 ( .A(TDSTARTADR[21]), .B(CACHE_ADDR1[16]), .Y(n2384) );
    zxo2b U765 ( .A(TDSTARTADR[18]), .B(CACHE_ADDR1[13]), .Y(n2388) );
    zxo2b U766 ( .A(TDSTARTADR[19]), .B(CACHE_ADDR1[14]), .Y(n2387) );
    zxo2b U767 ( .A(TDSTARTADR[16]), .B(CACHE_ADDR1[11]), .Y(n2390) );
    zxo2b U768 ( .A(TDSTARTADR[17]), .B(CACHE_ADDR1[12]), .Y(n2389) );
    zxo2b U769 ( .A(n2175), .B(TDSTARTADR[25]), .Y(n2415) );
    zxo2b U770 ( .A(n2174), .B(TDSTARTADR[22]), .Y(n2416) );
    zxo2b U771 ( .A(n2173), .B(TDSTARTADR[19]), .Y(n2417) );
    zxo2b U772 ( .A(n2178), .B(TDSTARTADR[31]), .Y(n2428) );
    zxo2b U773 ( .A(n2176), .B(TDSTARTADR[14]), .Y(n2427) );
    zxo2b U774 ( .A(n2177), .B(TDSTARTADR[21]), .Y(n2426) );
    zxo2b U775 ( .A(n2185), .B(TDSTARTADR[23]), .Y(n2419) );
    zxo2b U776 ( .A(n2183), .B(TDSTARTADR[6]), .Y(n2420) );
    zxo2b U777 ( .A(n2181), .B(TDSTARTADR[5]), .Y(n2421) );
    zxo2b U778 ( .A(n2179), .B(TDSTARTADR[7]), .Y(n2422) );
    zxo2b U779 ( .A(n2188), .B(TDSTARTADR[8]), .Y(n2425) );
    zxo2b U780 ( .A(n2186), .B(TDSTARTADR[15]), .Y(n2424) );
    zxo2b U781 ( .A(n2187), .B(TDSTARTADR[20]), .Y(n2423) );
    zxo2b U782 ( .A(CACHE_ADDR2[24]), .B(TDSTARTADR[29]), .Y(n2371) );
    zxo2b U783 ( .A(CACHE_ADDR2[23]), .B(TDSTARTADR[28]), .Y(n2372) );
    zxo2b U784 ( .A(CACHE_ADDR2[21]), .B(TDSTARTADR[26]), .Y(n2369) );
    zxo2b U785 ( .A(CACHE_ADDR2[25]), .B(TDSTARTADR[30]), .Y(n2370) );
    zxo2b U786 ( .A(CACHE_ADDR2[22]), .B(TDSTARTADR[27]), .Y(n2375) );
    zxo2b U787 ( .A(CACHE_ADDR2[13]), .B(TDSTARTADR[18]), .Y(n2374) );
    zxo2b U788 ( .A(CACHE_ADDR2[19]), .B(TDSTARTADR[24]), .Y(n2373) );
    zxo2b U789 ( .A(CACHE_ADDR2[11]), .B(TDSTARTADR[16]), .Y(n2377) );
    zxo2b U790 ( .A(CACHE_ADDR2[12]), .B(TDSTARTADR[17]), .Y(n2376) );
    zxo2b U791 ( .A(CACHE_ADDR2[7]), .B(TDSTARTADR[12]), .Y(n2379) );
    zxo2b U792 ( .A(CACHE_ADDR2[8]), .B(TDSTARTADR[13]), .Y(n2378) );
    zxo2b U793 ( .A(PHCI_DW1[0]), .B(RECOVERYMODE), .Y(n2391) );
    zor2b U794 ( .A(PERIOD_EN), .B(n2199), .Y(n2468) );
    zan2b U795 ( .A(TDIDLE1), .B(n2164), .Y(n2163) );
    zan2b U796 ( .A(TDIDLE2), .B(n2162), .Y(n2161) );
    zxo2b U797 ( .A(TDSTARTADR[11]), .B(CACHE_ADDR1[6]), .Y(n2220) );
    zxo2b U798 ( .A(TDSTARTADR[7]), .B(CACHE_ADDR1[2]), .Y(n2221) );
    zxo2b U799 ( .A(TDSTARTADR[12]), .B(CACHE_ADDR1[7]), .Y(n2222) );
    znd8b U800 ( .A(n2439), .B(n2440), .C(n2441), .D(n2434), .E(n2442), .F(
        n2443), .G(n2444), .H(n2430), .Y(n2225) );
    zxo2b U801 ( .A(CACHE_ADDR2[5]), .B(TDSTARTADR[10]), .Y(n2201) );
    zxo2b U802 ( .A(CACHE_ADDR2[4]), .B(TDSTARTADR[9]), .Y(n2202) );
    zxo2b U803 ( .A(CACHE_ADDR2[6]), .B(TDSTARTADR[11]), .Y(n2203) );
    znd8b U804 ( .A(n2423), .B(n2424), .C(n2425), .D(n2418), .E(n2426), .F(
        n2427), .G(n2428), .H(n2414), .Y(n2206) );
    zan2b U805 ( .A(n2146), .B(TDIDLE1), .Y(n2145) );
    zor2b U806 ( .A(n2151), .B(n2153), .Y(n2349) );
    zmux21lb U807 ( .A(n2133), .B(n2132), .S(TD_ACT2), .Y(n2397) );
    zxo2b U808 ( .A(n2335), .B(FRNUM_PER[3]), .Y(n2453) );
    zivb U809 ( .A(FRNUM[3]), .Y(n2335) );
    zxo2b U810 ( .A(n2334), .B(FRNUM_PER[4]), .Y(n2454) );
    zivb U811 ( .A(FRNUM[4]), .Y(n2334) );
    zxo2b U812 ( .A(n2333), .B(FRNUM_PER[6]), .Y(n2455) );
    zivb U813 ( .A(FRNUM[6]), .Y(n2333) );
    zxo2b U814 ( .A(n2331), .B(FRNUM_PER[7]), .Y(n2456) );
    zivb U815 ( .A(FRNUM[7]), .Y(n2331) );
    zxo2b U816 ( .A(n2338), .B(FRNUM_PER[1]), .Y(n2459) );
    zivb U817 ( .A(FRNUM[1]), .Y(n2338) );
    zxo2b U818 ( .A(n2336), .B(FRNUM[0]), .Y(n2458) );
    zxo2b U819 ( .A(n2337), .B(FRNUM[2]), .Y(n2457) );
    zor2b U820 ( .A(n2246), .B(n2247), .Y(n2248) );
    zivb U821 ( .A(n2246), .Y(n2467) );
    zor2b U822 ( .A(n2244), .B(n2391), .Y(n2469) );
    zan3b U823 ( .A(n2128), .B(n2129), .C(n2130), .Y(n2127) );
    zor2b U824 ( .A(n2022), .B(n2027), .Y(n2130) );
    zivb U825 ( .A(n2130), .Y(n2255) );
    zivb U826 ( .A(PARSETDEND2), .Y(n2129) );
    zivb U827 ( .A(PARSETDEND1), .Y(n2128) );
    zao33b U828 ( .A(TDIDLE1), .B(CACHEHIT1), .C(n2232), .D(TDIDLE2), .E(
        CACHEHIT2), .F(n2468), .Y(n2123) );
    zivb U829 ( .A(n2247), .Y(LAT_SAVEPLACE_COND) );
    zor2b U830 ( .A(FRNUM_PER[2]), .B(FRNUM_PER[1]), .Y(n2244) );
    zivb U831 ( .A(PHCI_DW1[0]), .Y(n2250) );
    zan2b U832 ( .A(n2015), .B(n2121), .Y(n2158) );
    zor2b U833 ( .A(PHASE_ParseTD), .B(PERIOD_END), .Y(n2170) );
    zxo2b U834 ( .A(n2168), .B(n2169), .Y(n2167) );
    zao21b U835 ( .A(TDSTARTADR[0]), .B(TDIDLE2), .C(n2146), .Y(n2160) );
    zivb U836 ( .A(n2232), .Y(n2146) );
    zor2b U837 ( .A(PERIOD_EN), .B(n2200), .Y(n2232) );
    zan2b U838 ( .A(n2140), .B(n2141), .Y(n2139) );
    zor2b U839 ( .A(FETCHTD), .B(PERIODSM_5), .Y(n2171) );
    zivb U840 ( .A(n2171), .Y(n2169) );
    zmux21lb U841 ( .A(n2161), .B(n2163), .S(CACHE_SEL), .Y(n2394) );
    zmux21lb U842 ( .A(PERIOD_EN), .B(PERIOD_RUN), .S(n2136), .Y(n2398) );
    zan2b U843 ( .A(n2137), .B(n2138), .Y(n2136) );
    zor2b U844 ( .A(CACHEHIT2), .B(CACHEHIT1), .Y(CACHE_HIT) );
    zivb U845 ( .A(n2164), .Y(CACHEHIT2) );
    zivb U846 ( .A(n2162), .Y(CACHEHIT1) );
    zor2b U847 ( .A(TDSTARTADR[0]), .B(n2025), .Y(n2226) );
    zmux21lb U848 ( .A(TDIDLE2), .B(n2232), .S(TDIDLE1), .Y(n2393) );
    zivb U849 ( .A(CACHE_HIT), .Y(n2152) );
    zivb U850 ( .A(n2237), .Y(n2447) );
    zor2b U851 ( .A(n2027), .B(n2144), .Y(n2237) );
    zivb U852 ( .A(n2230), .Y(n2446) );
    zmux21lb U853 ( .A(n2395), .B(n2396), .S(TD_ACT2), .Y(n2125) );
    zor2b U854 ( .A(TDPARSING1), .B(n2242), .Y(n2395) );
    zivb U855 ( .A(TDPARSING2), .Y(n2242) );
    zor2b U856 ( .A(TDPARSING2), .B(n2243), .Y(n2396) );
    zivb U857 ( .A(TDPARSING1), .Y(n2243) );
    zor2b U858 ( .A(TDHCIREQ1), .B(TDHCIREQ2), .Y(n2159) );
    zor2b U859 ( .A(PERIODSM_6), .B(n2170), .Y(n2168) );
    zan2b U860 ( .A(n2015), .B(n2121), .Y(n2154) );
    zivb U861 ( .A(n2226), .Y(n2122) );
    zor2b U862 ( .A(n2235), .B(n2236), .Y(n2155) );
    zxo2b U863 ( .A(FRLSTSIZE[1]), .B(FRLSTSIZE[0]), .Y(n2392) );
    zor2b U864 ( .A(n2165), .B(n2238), .Y(n2240) );
    zor2b U865 ( .A(CACHE_SEL_PRE), .B(n2238), .Y(n2241) );
    zivb U866 ( .A(n2413), .Y(n2470) );
    zxo2b U867 ( .A(TD_ACT1), .B(n2397), .Y(n2413) );
    znd8b U868 ( .A(n2340), .B(n2341), .C(n2342), .D(n2343), .E(n2344), .F(
        n2345), .G(n2346), .H(n2347), .Y(n2339) );
    zxo2b U869 ( .A(n2327), .B(FRNUM_PER[10]), .Y(n2340) );
    zivb U870 ( .A(FRNUM[10]), .Y(n2327) );
    zxo2b U871 ( .A(n2325), .B(FRNUM_PER[8]), .Y(n2341) );
    zivb U872 ( .A(FRNUM[8]), .Y(n2325) );
    zxo2b U873 ( .A(n2329), .B(FRNUM_PER[9]), .Y(n2342) );
    zivb U874 ( .A(FRNUM[9]), .Y(n2329) );
    zxo2b U875 ( .A(n2323), .B(FRNUM_PER[11]), .Y(n2343) );
    zivb U876 ( .A(FRNUM[11]), .Y(n2323) );
    zxo2b U877 ( .A(n2319), .B(FRNUM_PER[5]), .Y(n2344) );
    zivb U878 ( .A(FRNUM[5]), .Y(n2319) );
    zivb U879 ( .A(FRNUM[13]), .Y(n2345) );
    zxo2b U880 ( .A(n2321), .B(FRNUM_PER[12]), .Y(n2346) );
    zivb U881 ( .A(FRNUM[12]), .Y(n2321) );
    zxo2b add_250_U1_1_12 ( .A(FRNUM[12]), .B(add_250_carry_12), .Y(
        FRNUM_PER_PRE574_12) );
    zhadrb add_250_U1_1_11 ( .A(FRNUM[11]), .B(add_250_carry_11), .CO(
        add_250_carry_12), .S(FRNUM_PER_PRE574_11) );
    zhadrb add_250_U1_1_10 ( .A(FRNUM[10]), .B(add_250_carry_10), .CO(
        add_250_carry_11), .S(FRNUM_PER_PRE574_10) );
    zhadrb add_250_U1_1_9 ( .A(FRNUM[9]), .B(add_250_carry_9), .CO(
        add_250_carry_10), .S(FRNUM_PER_PRE574_9) );
    zhadrb add_250_U1_1_8 ( .A(FRNUM[8]), .B(add_250_carry_8), .CO(
        add_250_carry_9), .S(FRNUM_PER_PRE574_8) );
    zhadrb add_250_U1_1_7 ( .A(FRNUM[7]), .B(add_250_carry_7), .CO(
        add_250_carry_8), .S(FRNUM_PER_PRE574_7) );
    zhadrb add_250_U1_1_6 ( .A(FRNUM[6]), .B(add_250_carry_6), .CO(
        add_250_carry_7), .S(FRNUM_PER_PRE574_6) );
    zhadrb add_250_U1_1_5 ( .A(FRNUM[5]), .B(add_250_carry_5), .CO(
        add_250_carry_6), .S(FRNUM_PER_PRE574_5) );
    zhadrb add_250_U1_1_4 ( .A(FRNUM[4]), .B(add_250_carry_4), .CO(
        add_250_carry_5), .S(FRNUM_PER_PRE574_4) );
    zhadrb add_250_U1_1_3 ( .A(FRNUM[3]), .B(add_250_carry_3), .CO(
        add_250_carry_4), .S(FRNUM_PER_PRE574_3) );
    zhadrb add_250_U1_1_2 ( .A(FRNUM[2]), .B(add_250_carry_2), .CO(
        add_250_carry_3), .S(FRNUM_PER_PRE574_2) );
    zhadrb add_250_U1_1_1 ( .A(FRNUM[1]), .B(FRNUM[0]), .CO(add_250_carry_2), 
        .S(FRNUM_PER_PRE574_1) );
    zivc U882 ( .A(n2355), .Y(n2118) );
    zor2b U883 ( .A(n2356), .B(n2117), .Y(n2355) );
    zivb U884 ( .A(n2352), .Y(n2356) );
    zivb U885 ( .A(FRNUM[0]), .Y(FRNUM_PER_PRE574_0) );
    zivc U886 ( .A(n2354), .Y(n2119) );
    zor2b U887 ( .A(n2352), .B(n2117), .Y(n2354) );
    zmux21lb U888 ( .A(n2267), .B(n2268), .S(n2033), .Y(SAVEPTR679_31) );
    zivb U889 ( .A(PHCI_DW0[31]), .Y(n2268) );
    zmux21lb U890 ( .A(n2269), .B(n2270), .S(n2033), .Y(SAVEPTR679_30) );
    zivb U891 ( .A(PHCI_DW0[30]), .Y(n2270) );
    zmux21lb U892 ( .A(n2273), .B(n2274), .S(n2474), .Y(SAVEPTR679_29) );
    zivb U893 ( .A(PHCI_DW0[29]), .Y(n2274) );
    zmux21lb U894 ( .A(n2275), .B(n2276), .S(n2475), .Y(SAVEPTR679_28) );
    zivb U895 ( .A(PHCI_DW0[28]), .Y(n2276) );
    zmux21lb U896 ( .A(n2277), .B(n2278), .S(n2033), .Y(SAVEPTR679_27) );
    zivb U897 ( .A(PHCI_DW0[27]), .Y(n2278) );
    zmux21lb U898 ( .A(n2279), .B(n2280), .S(n2033), .Y(SAVEPTR679_26) );
    zivb U899 ( .A(PHCI_DW0[26]), .Y(n2280) );
    zmux21lb U900 ( .A(n2281), .B(n2282), .S(n2473), .Y(SAVEPTR679_25) );
    zivb U901 ( .A(PHCI_DW0[25]), .Y(n2282) );
    zmux21lb U902 ( .A(n2283), .B(n2284), .S(n2474), .Y(SAVEPTR679_24) );
    zivb U903 ( .A(PHCI_DW0[24]), .Y(n2284) );
    zmux21lb U904 ( .A(n2285), .B(n2286), .S(n2475), .Y(SAVEPTR679_23) );
    zivb U905 ( .A(PHCI_DW0[23]), .Y(n2286) );
    zmux21lb U906 ( .A(n2287), .B(n2288), .S(n2033), .Y(SAVEPTR679_22) );
    zivb U907 ( .A(PHCI_DW0[22]), .Y(n2288) );
    zmux21lb U908 ( .A(n2289), .B(n2290), .S(n2033), .Y(SAVEPTR679_21) );
    zivb U909 ( .A(PHCI_DW0[21]), .Y(n2290) );
    zmux21lb U910 ( .A(n2291), .B(n2292), .S(n2473), .Y(SAVEPTR679_20) );
    zivb U911 ( .A(PHCI_DW0[20]), .Y(n2292) );
    zmux21lb U912 ( .A(n2294), .B(n2295), .S(n2475), .Y(SAVEPTR679_19) );
    zivb U913 ( .A(PHCI_DW0[19]), .Y(n2295) );
    zmux21lb U914 ( .A(n2296), .B(n2297), .S(n2033), .Y(SAVEPTR679_18) );
    zivb U915 ( .A(PHCI_DW0[18]), .Y(n2297) );
    zmux21lb U916 ( .A(n2298), .B(n2299), .S(n2033), .Y(SAVEPTR679_17) );
    zivb U917 ( .A(PHCI_DW0[17]), .Y(n2299) );
    zmux21lb U918 ( .A(n2300), .B(n2301), .S(n2473), .Y(SAVEPTR679_16) );
    zivb U919 ( .A(PHCI_DW0[16]), .Y(n2301) );
    zmux21lb U920 ( .A(n2302), .B(n2303), .S(n2474), .Y(SAVEPTR679_15) );
    zivb U921 ( .A(PHCI_DW0[15]), .Y(n2303) );
    zmux21lb U922 ( .A(n2304), .B(n2305), .S(n2475), .Y(SAVEPTR679_14) );
    zivb U923 ( .A(PHCI_DW0[14]), .Y(n2305) );
    zmux21lb U924 ( .A(n2306), .B(n2307), .S(n2033), .Y(SAVEPTR679_13) );
    zivb U925 ( .A(PHCI_DW0[13]), .Y(n2307) );
    zmux21lb U926 ( .A(n2308), .B(n2309), .S(n2033), .Y(SAVEPTR679_12) );
    zivb U927 ( .A(PHCI_DW0[12]), .Y(n2309) );
    zmux21lb U928 ( .A(n2310), .B(n2311), .S(n2473), .Y(SAVEPTR679_11) );
    zivb U929 ( .A(PHCI_DW0[11]), .Y(n2311) );
    zmux21lb U930 ( .A(n2312), .B(n2313), .S(n2474), .Y(SAVEPTR679_10) );
    zivb U931 ( .A(PHCI_DW0[10]), .Y(n2313) );
    zmux21lb U932 ( .A(n2252), .B(n2253), .S(n2475), .Y(SAVEPTR679_9) );
    zivb U933 ( .A(PHCI_DW0[9]), .Y(n2253) );
    zmux21lb U934 ( .A(n2257), .B(n2258), .S(n2033), .Y(SAVEPTR679_8) );
    zivb U935 ( .A(PHCI_DW0[8]), .Y(n2258) );
    zmux21lb U936 ( .A(n2259), .B(n2260), .S(n2033), .Y(SAVEPTR679_7) );
    zivb U937 ( .A(PHCI_DW0[7]), .Y(n2260) );
    zmux21lb U938 ( .A(n2261), .B(n2262), .S(n2473), .Y(SAVEPTR679_6) );
    zivb U939 ( .A(PHCI_DW0[6]), .Y(n2262) );
    zmux21lb U940 ( .A(n2263), .B(n2264), .S(n2474), .Y(SAVEPTR679_5) );
    zivb U941 ( .A(PHCI_DW0[5]), .Y(n2264) );
    zmux21lb U942 ( .A(n2265), .B(n2266), .S(n2475), .Y(SAVEPTR679_4) );
    zivb U943 ( .A(PHCI_DW0[4]), .Y(n2266) );
    zmux21lb U944 ( .A(n2271), .B(n2272), .S(n2473), .Y(SAVEPTR679_3) );
    zivb U945 ( .A(PHCI_DW0[3]), .Y(n2272) );
    zbfb U946 ( .A(n2033), .Y(n2473) );
    zmux21lb U947 ( .A(n2293), .B(n2236), .S(n2474), .Y(SAVEPTR679_2) );
    zivb U948 ( .A(PHCI_DW0[2]), .Y(n2236) );
    zmux21lb U949 ( .A(n2314), .B(n2235), .S(n2475), .Y(SAVEPTR679_1) );
    zivb U950 ( .A(PHCI_DW0[1]), .Y(n2235) );
    zbfb U951 ( .A(n2033), .Y(n2475) );
    zmux21lb U952 ( .A(n2315), .B(n2316), .S(n2033), .Y(SAVEPTR679_0) );
    zivb U953 ( .A(PHCI_DW0[0]), .Y(n2316) );
    zor2b U954 ( .A(n2099), .B(n2100), .Y(TDSTARTADR717_31) );
    zor2b U955 ( .A(n2097), .B(n2098), .Y(TDSTARTADR717_30) );
    zor2b U956 ( .A(n2095), .B(n2096), .Y(TDSTARTADR717_29) );
    zor2b U957 ( .A(n2093), .B(n2094), .Y(TDSTARTADR717_28) );
    zor2b U958 ( .A(n2091), .B(n2092), .Y(TDSTARTADR717_27) );
    zor2b U959 ( .A(n2089), .B(n2090), .Y(TDSTARTADR717_26) );
    zor2b U960 ( .A(n2087), .B(n2088), .Y(TDSTARTADR717_25) );
    zor2b U961 ( .A(n2085), .B(n2086), .Y(TDSTARTADR717_24) );
    zor2b U962 ( .A(n2083), .B(n2084), .Y(TDSTARTADR717_23) );
    zor2b U963 ( .A(n2081), .B(n2082), .Y(TDSTARTADR717_22) );
    zor2b U964 ( .A(n2079), .B(n2080), .Y(TDSTARTADR717_21) );
    zor2b U965 ( .A(n2077), .B(n2078), .Y(TDSTARTADR717_20) );
    zor2b U966 ( .A(n2075), .B(n2076), .Y(TDSTARTADR717_19) );
    zor2b U967 ( .A(n2073), .B(n2074), .Y(TDSTARTADR717_18) );
    zor2b U968 ( .A(n2071), .B(n2072), .Y(TDSTARTADR717_17) );
    zor2b U969 ( .A(n2069), .B(n2070), .Y(TDSTARTADR717_16) );
    zor2b U970 ( .A(n2067), .B(n2068), .Y(TDSTARTADR717_15) );
    zor2b U971 ( .A(n2065), .B(n2066), .Y(TDSTARTADR717_14) );
    zor2b U972 ( .A(n2063), .B(n2064), .Y(TDSTARTADR717_13) );
    zor2b U973 ( .A(n2061), .B(n2062), .Y(TDSTARTADR717_12) );
    zor2b U974 ( .A(n2059), .B(n2060), .Y(TDSTARTADR717_11) );
    zor2b U975 ( .A(n2057), .B(n2058), .Y(TDSTARTADR717_10) );
    zor2b U976 ( .A(n2055), .B(n2056), .Y(TDSTARTADR717_9) );
    zor2b U977 ( .A(n2053), .B(n2054), .Y(TDSTARTADR717_8) );
    zor2b U978 ( .A(n2051), .B(n2052), .Y(TDSTARTADR717_7) );
    zor2b U979 ( .A(n2049), .B(n2050), .Y(TDSTARTADR717_6) );
    zor2b U980 ( .A(n2047), .B(n2048), .Y(TDSTARTADR717_5) );
    zor2b U981 ( .A(n2045), .B(n2046), .Y(TDSTARTADR717_4) );
    zor2b U982 ( .A(n2043), .B(n2044), .Y(TDSTARTADR717_3) );
    zor2b U983 ( .A(n2041), .B(n2042), .Y(TDSTARTADR717_2) );
    zivd U984 ( .A(n2248), .Y(n2483) );
    zivd U985 ( .A(n2256), .Y(n2131) );
    zor2b U986 ( .A(n2039), .B(n2040), .Y(TDSTARTADR717_1) );
    zivd U987 ( .A(n2251), .Y(n2448) );
    zivd U988 ( .A(n2248), .Y(n2449) );
    zivd U989 ( .A(n2254), .Y(n2451) );
    zan2b U990 ( .A(DW1_0[0]), .B(n2478), .Y(n2037) );
    zivd U991 ( .A(n2256), .Y(n2478) );
    zivd U992 ( .A(n2254), .Y(n2479) );
    zivd U993 ( .A(n2251), .Y(n2480) );
    zivb U994 ( .A(n2367), .Y(n2366) );
    zivb U995 ( .A(n2363), .Y(n2362) );
    zao22b U996 ( .A(FROZEN), .B(n2025), .C(n2028), .D(n2029), .Y(FROZEN1654)
         );
    zmux21lb U997 ( .A(n2199), .B(n2200), .S(TD_ACT2), .Y(n2028) );
    zivb U998 ( .A(n2126), .Y(n2029) );
    zor2b U999 ( .A(RUN), .B(n2137), .Y(n2126) );
    zmux21lb U1000 ( .A(n2409), .B(n2410), .S(ITDIDLE2), .Y(EXEITD21109) );
    zivb U1001 ( .A(n2238), .Y(PHASENXT_ParseTD) );
    zoai21b U1002 ( .A(n2120), .B(n2239), .C(n2109), .Y(n2238) );
    zor2b U1003 ( .A(n2032), .B(n2474), .Y(RECOVERYMODE642) );
    zmux21lb U1004 ( .A(n2405), .B(n2406), .S(QHIDLE2), .Y(EXEQH21183) );
    zao22b U1005 ( .A(PHASENXT_FetchTD), .B(n2115), .C(DWNUM[2]), .D(n2112), 
        .Y(DWNUM1434_2) );
    zao22b U1006 ( .A(PHASENXT_FetchTD), .B(n2116), .C(DWNUM[3]), .D(n2112), 
        .Y(DWNUM1434_3) );
    zmux21lb U1007 ( .A(n2403), .B(n2404), .S(SITDIDLE1), .Y(EXESITD11220) );
    zor2b U1008 ( .A(TDCMDSTART1), .B(TDCMDSTART2), .Y(TRANEXED1556) );
    zivb U1009 ( .A(n2143), .Y(n2103) );
    zan3b U1010 ( .A(TDIDLE1), .B(n2121), .C(n2160), .Y(n2105) );
    zivb U1011 ( .A(n2227), .Y(n2121) );
    zivb U1012 ( .A(n2165), .Y(CACHE_SEL_PRE) );
    zxo2b U1013 ( .A(n2166), .B(CACHE_SEL), .Y(n2165) );
    zmux21lb U1014 ( .A(n2407), .B(n2408), .S(QHIDLE1), .Y(EXEQH11146) );
    zivb U1015 ( .A(n2141), .Y(PERIOD_RUN_pre) );
    zor2b U1016 ( .A(n2025), .B(n2398), .Y(n2141) );
    zmux21lb U1017 ( .A(n2411), .B(n2412), .S(ITDIDLE1), .Y(EXEITD11072) );
    zao22b U1018 ( .A(PHASENXT_FetchTD), .B(n2114), .C(DWNUM[1]), .D(n2112), 
        .Y(DWNUM1434_1) );
    zao21b U1019 ( .A(n2359), .B(n2360), .C(n2231), .Y(n2358) );
    zor2b U1020 ( .A(n2116), .B(n2115), .Y(n2114) );
    zivb U1021 ( .A(n2114), .Y(n2348) );
    zivb U1022 ( .A(RUN), .Y(n2025) );
    zmux21lb U1023 ( .A(n2401), .B(n2402), .S(SITDIDLE2), .Y(EXESITD21257) );
    zxo2b U1024 ( .A(TD_ACT2), .B(n2124), .Y(TD_ACT_SEL827) );
    zan2b U1025 ( .A(n2125), .B(n2126), .Y(n2124) );
    zivb U1026 ( .A(FETCHTDNXT), .Y(n2112) );
    zivb U1027 ( .A(n2358), .Y(PHASENXT_FetchTD) );
    zivb U1028 ( .A(n2148), .Y(n2156) );
    zivb U1029 ( .A(n2159), .Y(n2157) );
    zivb U1030 ( .A(n2231), .Y(n2109) );
    zao21b U1031 ( .A(EXE_HALT), .B(n2137), .C(GEN_PERR), .Y(n2231) );
    zivb U1032 ( .A(SWDBG), .Y(n2137) );
    zan2b U1033 ( .A(n2034), .B(n2035), .Y(FRNUM_INC506) );
    zivb U1034 ( .A(LIST_SEL), .Y(n2351) );
    zor2b U1035 ( .A(PERIOD_ACT), .B(PERIOD_RUN), .Y(n2035) );
    zivb U1036 ( .A(n2035), .Y(n2353) );
    zivb U1037 ( .A(n2200), .Y(TDIDLE2) );
    zivb U1038 ( .A(SITDIDLE2), .Y(n2193) );
    zivb U1039 ( .A(QHIDLE2), .Y(n2194) );
    zivb U1040 ( .A(ITDIDLE2), .Y(n2195) );
    zivc U1041 ( .A(n2199), .Y(TDIDLE1) );
    zivb U1042 ( .A(SITDIDLE1), .Y(n2196) );
    zivb U1043 ( .A(QHIDLE1), .Y(n2197) );
    zivb U1044 ( .A(ITDIDLE1), .Y(n2198) );
    zao21b U1045 ( .A(TRANEXED), .B(SWDBG), .C(GEN_PERR), .Y(RUN_C) );
    zan2b U1046 ( .A(CACHE_SEL), .B(n2022), .Y(CACHE_EN2) );
    zan2b U1047 ( .A(n2023), .B(n2022), .Y(CACHE_EN1) );
    zan2b U1048 ( .A(n2472), .B(FRNUM_PER[3]), .Y(PERHCIADR[2]) );
    zan2b U1049 ( .A(PHASENXT_FetchPList), .B(FRNUM_PER[4]), .Y(PERHCIADR[3])
         );
    zan2b U1050 ( .A(n2472), .B(FRNUM_PER[5]), .Y(PERHCIADR[4]) );
    zmux21lb U1051 ( .A(n2182), .B(n2332), .S(n2472), .Y(PERHCIADR[5]) );
    zmux21lb U1052 ( .A(n2184), .B(n2330), .S(PHASENXT_FetchPList), .Y(
        PERHCIADR[6]) );
    zmux21lb U1053 ( .A(n2180), .B(n2324), .S(n2472), .Y(PERHCIADR[7]) );
    zmux21lb U1054 ( .A(n2189), .B(n2328), .S(PHASENXT_FetchPList), .Y(
        PERHCIADR[8]) );
    zmux21lb U1055 ( .A(n2191), .B(n2326), .S(n2472), .Y(PERHCIADR[9]) );
    zmux21lb U1056 ( .A(n2190), .B(n2400), .S(n2472), .Y(PERHCIADR[10]) );
    zao21b U1057 ( .A(FRLSTSIZE[1]), .B(n2462), .C(n2322), .Y(n2400) );
    zivb U1058 ( .A(FRLSTSIZE[0]), .Y(n2462) );
    zivb U1059 ( .A(n2400), .Y(FRNUM_PER[11]) );
    zmux21lb U1060 ( .A(n2192), .B(n2399), .S(PHASENXT_FetchPList), .Y(
        PERHCIADR[11]) );
    zor2b U1061 ( .A(n2320), .B(n2392), .Y(n2399) );
    zivb U1062 ( .A(n2399), .Y(FRNUM_PER[12]) );
    zmux21hb U1063 ( .A(TDSTARTADR[12]), .B(FLBASE[0]), .S(PHASENXT_FetchPList
        ), .Y(PERHCIADR[12]) );
    zmux21hb U1064 ( .A(TDSTARTADR[13]), .B(FLBASE[1]), .S(n2472), .Y(
        PERHCIADR[13]) );
    zmux21hb U1065 ( .A(TDSTARTADR[14]), .B(FLBASE[2]), .S(PHASENXT_FetchPList
        ), .Y(PERHCIADR[14]) );
    zmux21hb U1066 ( .A(TDSTARTADR[15]), .B(FLBASE[3]), .S(n2472), .Y(
        PERHCIADR[15]) );
    zmux21hb U1067 ( .A(TDSTARTADR[16]), .B(FLBASE[4]), .S(PHASENXT_FetchPList
        ), .Y(PERHCIADR[16]) );
    zmux21hb U1068 ( .A(TDSTARTADR[17]), .B(FLBASE[5]), .S(n2472), .Y(
        PERHCIADR[17]) );
    zmux21hb U1069 ( .A(TDSTARTADR[18]), .B(FLBASE[6]), .S(PHASENXT_FetchPList
        ), .Y(PERHCIADR[18]) );
    zmux21hb U1070 ( .A(TDSTARTADR[19]), .B(FLBASE[7]), .S(n2472), .Y(
        PERHCIADR[19]) );
    zmux21hb U1071 ( .A(TDSTARTADR[20]), .B(FLBASE[8]), .S(PHASENXT_FetchPList
        ), .Y(PERHCIADR[20]) );
    zmux21hb U1072 ( .A(TDSTARTADR[21]), .B(FLBASE[9]), .S(n2472), .Y(
        PERHCIADR[21]) );
    zmux21hb U1073 ( .A(TDSTARTADR[22]), .B(FLBASE[10]), .S(
        PHASENXT_FetchPList), .Y(PERHCIADR[22]) );
    zmux21hb U1074 ( .A(TDSTARTADR[23]), .B(FLBASE[11]), .S(n2472), .Y(
        PERHCIADR[23]) );
    zmux21hb U1075 ( .A(TDSTARTADR[24]), .B(FLBASE[12]), .S(
        PHASENXT_FetchPList), .Y(PERHCIADR[24]) );
    zmux21hb U1076 ( .A(TDSTARTADR[25]), .B(FLBASE[13]), .S(n2472), .Y(
        PERHCIADR[25]) );
    zmux21hb U1077 ( .A(TDSTARTADR[26]), .B(FLBASE[14]), .S(
        PHASENXT_FetchPList), .Y(PERHCIADR[26]) );
    zmux21hb U1078 ( .A(TDSTARTADR[27]), .B(FLBASE[15]), .S(n2472), .Y(
        PERHCIADR[27]) );
    zmux21hb U1079 ( .A(TDSTARTADR[28]), .B(FLBASE[16]), .S(
        PHASENXT_FetchPList), .Y(PERHCIADR[28]) );
    zmux21hb U1080 ( .A(TDSTARTADR[29]), .B(FLBASE[17]), .S(n2472), .Y(
        PERHCIADR[29]) );
    zmux21hb U1081 ( .A(TDSTARTADR[30]), .B(FLBASE[18]), .S(
        PHASENXT_FetchPList), .Y(PERHCIADR[30]) );
    zmux21hb U1082 ( .A(TDSTARTADR[31]), .B(FLBASE[19]), .S(n2472), .Y(
        PERHCIADR[31]) );
    zivd U1083 ( .A(n2350), .Y(n2472) );
    zor2b U1084 ( .A(n2142), .B(n2231), .Y(n2350) );
    zivd U1085 ( .A(n2350), .Y(PHASENXT_FetchPList) );
    zivb U1086 ( .A(n2463), .Y(TD_CACHE_EN2) );
    zor2b U1087 ( .A(n2228), .B(n2023), .Y(n2463) );
    zivb U1088 ( .A(n2465), .Y(TD_CACHE_EN1) );
    zor2b U1089 ( .A(CACHE_SEL), .B(n2228), .Y(n2465) );
    zan2b U1090 ( .A(n2021), .B(TD_ACT2), .Y(PER_EXE2) );
    zan2b U1091 ( .A(n2024), .B(TD_ACT1), .Y(PER_EXE1) );
    zor2b U1092 ( .A(PERIODSM_1), .B(PHASE_FetchFSTN), .Y(PCACHE_EN) );
    zivb U1093 ( .A(PCACHE_EN), .Y(n2022) );
    zor2b U1094 ( .A(n2011), .B(TD_PARSE_GO2_T), .Y(TD_PARSE_GO2) );
    zor2b U1095 ( .A(n2010), .B(TD_PARSE_GO1_T), .Y(TD_PARSE_GO1) );
    zor2b U1096 ( .A(PCACHE_EN), .B(PERIODSM_3), .Y(FETCHTD) );
    zivb U1097 ( .A(TDHCIREQ1), .Y(n2132) );
    zivb U1098 ( .A(TDHCIREQ2), .Y(n2133) );
    zivb U1099 ( .A(n2135), .Y(PHCI_PRESOF) );
    zdffqrb FRNUM_PER_PRE_reg_12 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_12), .R(
        TRST_), .Q(FRNUM_PER_PRE_12) );
    zivb U1100 ( .A(FRNUM_PER_PRE_12), .Y(n2320) );
    zdffqrb FRNUM_PER_PRE_reg_11 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_11), .R(
        TRST_), .Q(FRNUM_PER_PRE_11) );
    zivb U1101 ( .A(FRNUM_PER_PRE_11), .Y(n2322) );
    zdffqrb FRNUM_PER_PRE_reg_10 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_10), .R(
        TRST_), .Q(FRNUM_PER[10]) );
    zivb U1102 ( .A(FRNUM_PER[10]), .Y(n2326) );
    zdffqrb FRNUM_PER_PRE_reg_9 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_9), .R(
        TRST_), .Q(FRNUM_PER[9]) );
    zivb U1103 ( .A(FRNUM_PER[9]), .Y(n2328) );
    zdffqrb FRNUM_PER_PRE_reg_8 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_8), .R(
        TRST_), .Q(FRNUM_PER[8]) );
    zivb U1104 ( .A(FRNUM_PER[8]), .Y(n2324) );
    zdffqrb FRNUM_PER_PRE_reg_7 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_7), .R(
        TRST_), .Q(FRNUM_PER[7]) );
    zivb U1105 ( .A(FRNUM_PER[7]), .Y(n2330) );
    zdffqrb FRNUM_PER_PRE_reg_6 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_6), .R(
        TRST_), .Q(FRNUM_PER[6]) );
    zivb U1106 ( .A(FRNUM_PER[6]), .Y(n2332) );
    zdffqrb FRNUM_PER_PRE_reg_5 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_5), .R(
        TRST_), .Q(FRNUM_PER[5]) );
    zdffqrb FRNUM_PER_PRE_reg_4 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_4), .R(
        TRST_), .Q(FRNUM_PER[4]) );
    zdffqrb FRNUM_PER_PRE_reg_3 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_3), .R(
        TRST_), .Q(FRNUM_PER[3]) );
    zdffqrb FRNUM_PER_PRE_reg_2 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_2), .R(
        TRST_), .Q(FRNUM_PER[2]) );
    zivb U1107 ( .A(FRNUM_PER[2]), .Y(n2337) );
    zdffqrb FRNUM_PER_PRE_reg_1 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_1), .R(
        TRST_), .Q(FRNUM_PER[1]) );
    zdffqrb FRNUM_PER_PRE_reg_0 ( .CK(PCICLK), .D(FRNUM_PER_PRE597_0), .R(
        TRST_), .Q(FRNUM_PER[0]) );
    zivb U1108 ( .A(FRNUM_PER[0]), .Y(n2336) );
    zdffrb SAVEPTR_reg_31 ( .CK(PCICLK), .D(SAVEPTR679_31), .R(TRST_), .Q(
        SAVEPTR_31), .QN(n2267) );
    zdffrb SAVEPTR_reg_30 ( .CK(PCICLK), .D(SAVEPTR679_30), .R(TRST_), .Q(
        SAVEPTR_30), .QN(n2269) );
    zdffrb SAVEPTR_reg_29 ( .CK(PCICLK), .D(SAVEPTR679_29), .R(TRST_), .Q(
        SAVEPTR_29), .QN(n2273) );
    zdffrb SAVEPTR_reg_28 ( .CK(PCICLK), .D(SAVEPTR679_28), .R(TRST_), .Q(
        SAVEPTR_28), .QN(n2275) );
    zdffrb SAVEPTR_reg_27 ( .CK(PCICLK), .D(SAVEPTR679_27), .R(TRST_), .Q(
        SAVEPTR_27), .QN(n2277) );
    zdffrb SAVEPTR_reg_26 ( .CK(PCICLK), .D(SAVEPTR679_26), .R(TRST_), .Q(
        SAVEPTR_26), .QN(n2279) );
    zdffrb SAVEPTR_reg_25 ( .CK(PCICLK), .D(SAVEPTR679_25), .R(TRST_), .Q(
        SAVEPTR_25), .QN(n2281) );
    zdffrb SAVEPTR_reg_24 ( .CK(PCICLK), .D(SAVEPTR679_24), .R(TRST_), .Q(
        SAVEPTR_24), .QN(n2283) );
    zdffrb SAVEPTR_reg_23 ( .CK(PCICLK), .D(SAVEPTR679_23), .R(TRST_), .Q(
        SAVEPTR_23), .QN(n2285) );
    zdffrb SAVEPTR_reg_22 ( .CK(PCICLK), .D(SAVEPTR679_22), .R(TRST_), .Q(
        SAVEPTR_22), .QN(n2287) );
    zdffrb SAVEPTR_reg_21 ( .CK(PCICLK), .D(SAVEPTR679_21), .R(TRST_), .Q(
        SAVEPTR_21), .QN(n2289) );
    zdffrb SAVEPTR_reg_20 ( .CK(PCICLK), .D(SAVEPTR679_20), .R(TRST_), .Q(
        SAVEPTR_20), .QN(n2291) );
    zdffrb SAVEPTR_reg_19 ( .CK(PCICLK), .D(SAVEPTR679_19), .R(TRST_), .Q(
        SAVEPTR_19), .QN(n2294) );
    zdffrb SAVEPTR_reg_18 ( .CK(PCICLK), .D(SAVEPTR679_18), .R(TRST_), .Q(
        SAVEPTR_18), .QN(n2296) );
    zdffrb SAVEPTR_reg_17 ( .CK(PCICLK), .D(SAVEPTR679_17), .R(TRST_), .Q(
        SAVEPTR_17), .QN(n2298) );
    zdffrb SAVEPTR_reg_16 ( .CK(PCICLK), .D(SAVEPTR679_16), .R(TRST_), .Q(
        SAVEPTR_16), .QN(n2300) );
    zdffrb SAVEPTR_reg_15 ( .CK(PCICLK), .D(SAVEPTR679_15), .R(TRST_), .Q(
        SAVEPTR_15), .QN(n2302) );
    zdffrb SAVEPTR_reg_14 ( .CK(PCICLK), .D(SAVEPTR679_14), .R(TRST_), .Q(
        SAVEPTR_14), .QN(n2304) );
    zdffrb SAVEPTR_reg_13 ( .CK(PCICLK), .D(SAVEPTR679_13), .R(TRST_), .Q(
        SAVEPTR_13), .QN(n2306) );
    zdffrb SAVEPTR_reg_12 ( .CK(PCICLK), .D(SAVEPTR679_12), .R(TRST_), .Q(
        SAVEPTR_12), .QN(n2308) );
    zdffrb SAVEPTR_reg_11 ( .CK(PCICLK), .D(SAVEPTR679_11), .R(TRST_), .Q(
        SAVEPTR_11), .QN(n2310) );
    zdffrb SAVEPTR_reg_10 ( .CK(PCICLK), .D(SAVEPTR679_10), .R(TRST_), .Q(
        SAVEPTR_10), .QN(n2312) );
    zdffrb SAVEPTR_reg_9 ( .CK(PCICLK), .D(SAVEPTR679_9), .R(TRST_), .Q(
        SAVEPTR_9), .QN(n2252) );
    zdffrb SAVEPTR_reg_8 ( .CK(PCICLK), .D(SAVEPTR679_8), .R(TRST_), .Q(
        SAVEPTR_8), .QN(n2257) );
    zdffrb SAVEPTR_reg_7 ( .CK(PCICLK), .D(SAVEPTR679_7), .R(TRST_), .Q(
        SAVEPTR_7), .QN(n2259) );
    zdffrb SAVEPTR_reg_6 ( .CK(PCICLK), .D(SAVEPTR679_6), .R(TRST_), .Q(
        SAVEPTR_6), .QN(n2261) );
    zdffrb SAVEPTR_reg_5 ( .CK(PCICLK), .D(SAVEPTR679_5), .R(TRST_), .Q(
        SAVEPTR_5), .QN(n2263) );
    zdffrb SAVEPTR_reg_4 ( .CK(PCICLK), .D(SAVEPTR679_4), .R(TRST_), .Q(
        SAVEPTR_4), .QN(n2265) );
    zdffrb SAVEPTR_reg_3 ( .CK(PCICLK), .D(SAVEPTR679_3), .R(TRST_), .Q(
        SAVEPTR_3), .QN(n2271) );
    zdffrb SAVEPTR_reg_2 ( .CK(PCICLK), .D(SAVEPTR679_2), .R(TRST_), .Q(
        SAVEPTR_2), .QN(n2293) );
    zdffrb SAVEPTR_reg_1 ( .CK(PCICLK), .D(SAVEPTR679_1), .R(TRST_), .Q(
        SAVEPTR_1), .QN(n2314) );
    zdffrb SAVEPTR_reg_0 ( .CK(PCICLK), .D(SAVEPTR679_0), .R(TRST_), .Q(
        SAVEPTR_0), .QN(n2315) );
    zdffqrb TDSTARTADR_reg_31 ( .CK(PCICLK), .D(TDSTARTADR717_31), .R(TRST_), 
        .Q(TDSTARTADR[31]) );
    zdffqrb TDSTARTADR_reg_30 ( .CK(PCICLK), .D(TDSTARTADR717_30), .R(TRST_), 
        .Q(TDSTARTADR[30]) );
    zdffqrb TDSTARTADR_reg_29 ( .CK(PCICLK), .D(TDSTARTADR717_29), .R(TRST_), 
        .Q(TDSTARTADR[29]) );
    zdffqrb TDSTARTADR_reg_28 ( .CK(PCICLK), .D(TDSTARTADR717_28), .R(TRST_), 
        .Q(TDSTARTADR[28]) );
    zdffqrb TDSTARTADR_reg_27 ( .CK(PCICLK), .D(TDSTARTADR717_27), .R(TRST_), 
        .Q(TDSTARTADR[27]) );
    zdffqrb TDSTARTADR_reg_26 ( .CK(PCICLK), .D(TDSTARTADR717_26), .R(TRST_), 
        .Q(TDSTARTADR[26]) );
    zdffqrb TDSTARTADR_reg_25 ( .CK(PCICLK), .D(TDSTARTADR717_25), .R(TRST_), 
        .Q(TDSTARTADR[25]) );
    zdffqrb TDSTARTADR_reg_24 ( .CK(PCICLK), .D(TDSTARTADR717_24), .R(TRST_), 
        .Q(TDSTARTADR[24]) );
    zdffqrb TDSTARTADR_reg_23 ( .CK(PCICLK), .D(TDSTARTADR717_23), .R(TRST_), 
        .Q(TDSTARTADR[23]) );
    zdffqrb TDSTARTADR_reg_22 ( .CK(PCICLK), .D(TDSTARTADR717_22), .R(TRST_), 
        .Q(TDSTARTADR[22]) );
    zdffqrb TDSTARTADR_reg_21 ( .CK(PCICLK), .D(TDSTARTADR717_21), .R(TRST_), 
        .Q(TDSTARTADR[21]) );
    zdffqrb TDSTARTADR_reg_20 ( .CK(PCICLK), .D(TDSTARTADR717_20), .R(TRST_), 
        .Q(TDSTARTADR[20]) );
    zdffqrb TDSTARTADR_reg_19 ( .CK(PCICLK), .D(TDSTARTADR717_19), .R(TRST_), 
        .Q(TDSTARTADR[19]) );
    zdffqrb TDSTARTADR_reg_18 ( .CK(PCICLK), .D(TDSTARTADR717_18), .R(TRST_), 
        .Q(TDSTARTADR[18]) );
    zdffqrb TDSTARTADR_reg_17 ( .CK(PCICLK), .D(TDSTARTADR717_17), .R(TRST_), 
        .Q(TDSTARTADR[17]) );
    zdffqrb TDSTARTADR_reg_16 ( .CK(PCICLK), .D(TDSTARTADR717_16), .R(TRST_), 
        .Q(TDSTARTADR[16]) );
    zdffqrb TDSTARTADR_reg_15 ( .CK(PCICLK), .D(TDSTARTADR717_15), .R(TRST_), 
        .Q(TDSTARTADR[15]) );
    zdffqrb TDSTARTADR_reg_14 ( .CK(PCICLK), .D(TDSTARTADR717_14), .R(TRST_), 
        .Q(TDSTARTADR[14]) );
    zdffqrb TDSTARTADR_reg_13 ( .CK(PCICLK), .D(TDSTARTADR717_13), .R(TRST_), 
        .Q(TDSTARTADR[13]) );
    zdffqrb TDSTARTADR_reg_12 ( .CK(PCICLK), .D(TDSTARTADR717_12), .R(TRST_), 
        .Q(TDSTARTADR[12]) );
    zdffqrb TDSTARTADR_reg_11 ( .CK(PCICLK), .D(TDSTARTADR717_11), .R(TRST_), 
        .Q(TDSTARTADR[11]) );
    zivb U1109 ( .A(TDSTARTADR[11]), .Y(n2192) );
    zdffqrb TDSTARTADR_reg_10 ( .CK(PCICLK), .D(TDSTARTADR717_10), .R(TRST_), 
        .Q(TDSTARTADR[10]) );
    zivb U1110 ( .A(TDSTARTADR[10]), .Y(n2190) );
    zdffqrb TDSTARTADR_reg_9 ( .CK(PCICLK), .D(TDSTARTADR717_9), .R(TRST_), 
        .Q(TDSTARTADR[9]) );
    zivb U1111 ( .A(TDSTARTADR[9]), .Y(n2191) );
    zdffqrb TDSTARTADR_reg_8 ( .CK(PCICLK), .D(TDSTARTADR717_8), .R(TRST_), 
        .Q(TDSTARTADR[8]) );
    zivb U1112 ( .A(TDSTARTADR[8]), .Y(n2189) );
    zdffqrb TDSTARTADR_reg_7 ( .CK(PCICLK), .D(TDSTARTADR717_7), .R(TRST_), 
        .Q(TDSTARTADR[7]) );
    zivb U1113 ( .A(TDSTARTADR[7]), .Y(n2180) );
    zdffqrb TDSTARTADR_reg_6 ( .CK(PCICLK), .D(TDSTARTADR717_6), .R(TRST_), 
        .Q(TDSTARTADR[6]) );
    zivb U1114 ( .A(TDSTARTADR[6]), .Y(n2184) );
    zdffqrb TDSTARTADR_reg_5 ( .CK(PCICLK), .D(TDSTARTADR717_5), .R(TRST_), 
        .Q(TDSTARTADR[5]) );
    zivb U1115 ( .A(TDSTARTADR[5]), .Y(n2182) );
    zdffqrb TDSTARTADR_reg_4 ( .CK(PCICLK), .D(TDSTARTADR717_4), .R(TRST_), 
        .Q(TDSTARTADR[4]) );
    zdffqrb TDSTARTADR_reg_3 ( .CK(PCICLK), .D(TDSTARTADR717_3), .R(TRST_), 
        .Q(TDSTARTADR[3]) );
    zdffrb TDSTARTADR_reg_2 ( .CK(PCICLK), .D(TDSTARTADR717_2), .R(TRST_), .Q(
        TDSTARTADR[2]), .QN(n2116) );
    zdffqrb TDSTARTADR_reg_1 ( .CK(PCICLK), .D(TDSTARTADR717_1), .R(TRST_), 
        .Q(TDSTARTADR[1]) );
    zivb U1116 ( .A(TDSTARTADR[1]), .Y(n2115) );
    zdffqrb TDSTARTADR_reg_0 ( .CK(PCICLK), .D(TDSTARTADR717_0), .R(TRST_), 
        .Q(TDSTARTADR[0]) );
    zivb U1117 ( .A(TDSTARTADR[0]), .Y(n2317) );
    zdffqrb CACHE_ADDR1_reg_26 ( .CK(PCICLK), .D(CACHE_ADDR1996_26), .R(TRST_), 
        .Q(CACHE_ADDR1[26]) );
    zdffqrb CACHE_ADDR1_reg_25 ( .CK(PCICLK), .D(CACHE_ADDR1996_25), .R(TRST_), 
        .Q(CACHE_ADDR1[25]) );
    zivb U1118 ( .A(CACHE_ADDR1[25]), .Y(n2207) );
    zdffqrb CACHE_ADDR1_reg_24 ( .CK(PCICLK), .D(CACHE_ADDR1996_24), .R(TRST_), 
        .Q(CACHE_ADDR1[24]) );
    zivb U1119 ( .A(CACHE_ADDR1[24]), .Y(n2208) );
    zdffqrb CACHE_ADDR1_reg_23 ( .CK(PCICLK), .D(CACHE_ADDR1996_23), .R(TRST_), 
        .Q(CACHE_ADDR1[23]) );
    zivb U1120 ( .A(CACHE_ADDR1[23]), .Y(n2214) );
    zdffqrb CACHE_ADDR1_reg_22 ( .CK(PCICLK), .D(CACHE_ADDR1996_22), .R(TRST_), 
        .Q(CACHE_ADDR1[22]) );
    zdffqrb CACHE_ADDR1_reg_21 ( .CK(PCICLK), .D(CACHE_ADDR1996_21), .R(TRST_), 
        .Q(CACHE_ADDR1[21]) );
    zivb U1121 ( .A(CACHE_ADDR1[21]), .Y(n2216) );
    zdffqrb CACHE_ADDR1_reg_20 ( .CK(PCICLK), .D(CACHE_ADDR1996_20), .R(TRST_), 
        .Q(CACHE_ADDR1[20]) );
    zivb U1122 ( .A(CACHE_ADDR1[20]), .Y(n2219) );
    zdffqrb CACHE_ADDR1_reg_19 ( .CK(PCICLK), .D(CACHE_ADDR1996_19), .R(TRST_), 
        .Q(CACHE_ADDR1[19]) );
    zdffqrb CACHE_ADDR1_reg_18 ( .CK(PCICLK), .D(CACHE_ADDR1996_18), .R(TRST_), 
        .Q(CACHE_ADDR1[18]) );
    zdffqrb CACHE_ADDR1_reg_17 ( .CK(PCICLK), .D(CACHE_ADDR1996_17), .R(TRST_), 
        .Q(CACHE_ADDR1[17]) );
    zivb U1123 ( .A(CACHE_ADDR1[17]), .Y(n2212) );
    zdffqrb CACHE_ADDR1_reg_16 ( .CK(PCICLK), .D(CACHE_ADDR1996_16), .R(TRST_), 
        .Q(CACHE_ADDR1[16]) );
    zdffqrb CACHE_ADDR1_reg_15 ( .CK(PCICLK), .D(CACHE_ADDR1996_15), .R(TRST_), 
        .Q(CACHE_ADDR1[15]) );
    zivb U1124 ( .A(CACHE_ADDR1[15]), .Y(n2211) );
    zdffqrb CACHE_ADDR1_reg_14 ( .CK(PCICLK), .D(CACHE_ADDR1996_14), .R(TRST_), 
        .Q(CACHE_ADDR1[14]) );
    zdffqrb CACHE_ADDR1_reg_13 ( .CK(PCICLK), .D(CACHE_ADDR1996_13), .R(TRST_), 
        .Q(CACHE_ADDR1[13]) );
    zdffqrb CACHE_ADDR1_reg_12 ( .CK(PCICLK), .D(CACHE_ADDR1996_12), .R(TRST_), 
        .Q(CACHE_ADDR1[12]) );
    zdffqrb CACHE_ADDR1_reg_11 ( .CK(PCICLK), .D(CACHE_ADDR1996_11), .R(TRST_), 
        .Q(CACHE_ADDR1[11]) );
    zdffqrb CACHE_ADDR1_reg_10 ( .CK(PCICLK), .D(CACHE_ADDR1996_10), .R(TRST_), 
        .Q(CACHE_ADDR1[10]) );
    zdffqrb CACHE_ADDR1_reg_9 ( .CK(PCICLK), .D(CACHE_ADDR1996_9), .R(TRST_), 
        .Q(CACHE_ADDR1[9]) );
    zivb U1125 ( .A(CACHE_ADDR1[9]), .Y(n2210) );
    zdffqrb CACHE_ADDR1_reg_8 ( .CK(PCICLK), .D(CACHE_ADDR1996_8), .R(TRST_), 
        .Q(CACHE_ADDR1[8]) );
    zivb U1126 ( .A(CACHE_ADDR1[8]), .Y(n2213) );
    zdffqrb CACHE_ADDR1_reg_7 ( .CK(PCICLK), .D(CACHE_ADDR1996_7), .R(TRST_), 
        .Q(CACHE_ADDR1[7]) );
    zdffqrb CACHE_ADDR1_reg_6 ( .CK(PCICLK), .D(CACHE_ADDR1996_6), .R(TRST_), 
        .Q(CACHE_ADDR1[6]) );
    zdffqrb CACHE_ADDR1_reg_5 ( .CK(PCICLK), .D(CACHE_ADDR1996_5), .R(TRST_), 
        .Q(CACHE_ADDR1[5]) );
    zdffqrb CACHE_ADDR1_reg_4 ( .CK(PCICLK), .D(CACHE_ADDR1996_4), .R(TRST_), 
        .Q(CACHE_ADDR1[4]) );
    zivb U1127 ( .A(CACHE_ADDR1[4]), .Y(n2209) );
    zdffqrb CACHE_ADDR1_reg_3 ( .CK(PCICLK), .D(CACHE_ADDR1996_3), .R(TRST_), 
        .Q(CACHE_ADDR1[3]) );
    zivb U1128 ( .A(CACHE_ADDR1[3]), .Y(n2215) );
    zdffqrb CACHE_ADDR1_reg_2 ( .CK(PCICLK), .D(CACHE_ADDR1996_2), .R(TRST_), 
        .Q(CACHE_ADDR1[2]) );
    zdffqrb CACHE_ADDR1_reg_1 ( .CK(PCICLK), .D(CACHE_ADDR1996_1), .R(TRST_), 
        .Q(CACHE_ADDR1[1]) );
    zivb U1129 ( .A(CACHE_ADDR1[1]), .Y(n2218) );
    zdffqrb CACHE_ADDR1_reg_0 ( .CK(PCICLK), .D(CACHE_ADDR1996_0), .R(TRST_), 
        .Q(CACHE_ADDR1[0]) );
    zivb U1130 ( .A(CACHE_ADDR1[0]), .Y(n2217) );
    zdffqrb CACHE_ADDR2_reg_26 ( .CK(PCICLK), .D(CACHE_ADDR21034_26), .R(TRST_
        ), .Q(CACHE_ADDR2[26]) );
    zivb U1131 ( .A(CACHE_ADDR2[26]), .Y(n2178) );
    zdffqrb CACHE_ADDR2_reg_25 ( .CK(PCICLK), .D(CACHE_ADDR21034_25), .R(TRST_
        ), .Q(CACHE_ADDR2[25]) );
    zdffqrb CACHE_ADDR2_reg_24 ( .CK(PCICLK), .D(CACHE_ADDR21034_24), .R(TRST_
        ), .Q(CACHE_ADDR2[24]) );
    zdffqrb CACHE_ADDR2_reg_23 ( .CK(PCICLK), .D(CACHE_ADDR21034_23), .R(TRST_
        ), .Q(CACHE_ADDR2[23]) );
    zdffqrb CACHE_ADDR2_reg_22 ( .CK(PCICLK), .D(CACHE_ADDR21034_22), .R(TRST_
        ), .Q(CACHE_ADDR2[22]) );
    zdffqrb CACHE_ADDR2_reg_21 ( .CK(PCICLK), .D(CACHE_ADDR21034_21), .R(TRST_
        ), .Q(CACHE_ADDR2[21]) );
    zdffqrb CACHE_ADDR2_reg_20 ( .CK(PCICLK), .D(CACHE_ADDR21034_20), .R(TRST_
        ), .Q(CACHE_ADDR2[20]) );
    zivb U1132 ( .A(CACHE_ADDR2[20]), .Y(n2175) );
    zdffqrb CACHE_ADDR2_reg_19 ( .CK(PCICLK), .D(CACHE_ADDR21034_19), .R(TRST_
        ), .Q(CACHE_ADDR2[19]) );
    zdffqrb CACHE_ADDR2_reg_18 ( .CK(PCICLK), .D(CACHE_ADDR21034_18), .R(TRST_
        ), .Q(CACHE_ADDR2[18]) );
    zivb U1133 ( .A(CACHE_ADDR2[18]), .Y(n2185) );
    zdffqrb CACHE_ADDR2_reg_17 ( .CK(PCICLK), .D(CACHE_ADDR21034_17), .R(TRST_
        ), .Q(CACHE_ADDR2[17]) );
    zivb U1134 ( .A(CACHE_ADDR2[17]), .Y(n2174) );
    zdffqrb CACHE_ADDR2_reg_16 ( .CK(PCICLK), .D(CACHE_ADDR21034_16), .R(TRST_
        ), .Q(CACHE_ADDR2[16]) );
    zivb U1135 ( .A(CACHE_ADDR2[16]), .Y(n2177) );
    zdffqrb CACHE_ADDR2_reg_15 ( .CK(PCICLK), .D(CACHE_ADDR21034_15), .R(TRST_
        ), .Q(CACHE_ADDR2[15]) );
    zivb U1136 ( .A(CACHE_ADDR2[15]), .Y(n2187) );
    zdffqrb CACHE_ADDR2_reg_14 ( .CK(PCICLK), .D(CACHE_ADDR21034_14), .R(TRST_
        ), .Q(CACHE_ADDR2[14]) );
    zivb U1137 ( .A(CACHE_ADDR2[14]), .Y(n2173) );
    zdffqrb CACHE_ADDR2_reg_13 ( .CK(PCICLK), .D(CACHE_ADDR21034_13), .R(TRST_
        ), .Q(CACHE_ADDR2[13]) );
    zdffqrb CACHE_ADDR2_reg_12 ( .CK(PCICLK), .D(CACHE_ADDR21034_12), .R(TRST_
        ), .Q(CACHE_ADDR2[12]) );
    zdffqrb CACHE_ADDR2_reg_11 ( .CK(PCICLK), .D(CACHE_ADDR21034_11), .R(TRST_
        ), .Q(CACHE_ADDR2[11]) );
    zdffqrb CACHE_ADDR2_reg_10 ( .CK(PCICLK), .D(CACHE_ADDR21034_10), .R(TRST_
        ), .Q(CACHE_ADDR2[10]) );
    zivb U1138 ( .A(CACHE_ADDR2[10]), .Y(n2186) );
    zdffqrb CACHE_ADDR2_reg_9 ( .CK(PCICLK), .D(CACHE_ADDR21034_9), .R(TRST_), 
        .Q(CACHE_ADDR2[9]) );
    zivb U1139 ( .A(CACHE_ADDR2[9]), .Y(n2176) );
    zdffqrb CACHE_ADDR2_reg_8 ( .CK(PCICLK), .D(CACHE_ADDR21034_8), .R(TRST_), 
        .Q(CACHE_ADDR2[8]) );
    zdffqrb CACHE_ADDR2_reg_7 ( .CK(PCICLK), .D(CACHE_ADDR21034_7), .R(TRST_), 
        .Q(CACHE_ADDR2[7]) );
    zdffqrb CACHE_ADDR2_reg_6 ( .CK(PCICLK), .D(CACHE_ADDR21034_6), .R(TRST_), 
        .Q(CACHE_ADDR2[6]) );
    zdffqrb CACHE_ADDR2_reg_5 ( .CK(PCICLK), .D(CACHE_ADDR21034_5), .R(TRST_), 
        .Q(CACHE_ADDR2[5]) );
    zdffqrb CACHE_ADDR2_reg_4 ( .CK(PCICLK), .D(CACHE_ADDR21034_4), .R(TRST_), 
        .Q(CACHE_ADDR2[4]) );
    zdffqrb CACHE_ADDR2_reg_3 ( .CK(PCICLK), .D(CACHE_ADDR21034_3), .R(TRST_), 
        .Q(CACHE_ADDR2[3]) );
    zivb U1140 ( .A(CACHE_ADDR2[3]), .Y(n2188) );
    zdffqrb CACHE_ADDR2_reg_2 ( .CK(PCICLK), .D(CACHE_ADDR21034_2), .R(TRST_), 
        .Q(CACHE_ADDR2[2]) );
    zivb U1141 ( .A(CACHE_ADDR2[2]), .Y(n2179) );
    zdffqrb CACHE_ADDR2_reg_1 ( .CK(PCICLK), .D(CACHE_ADDR21034_1), .R(TRST_), 
        .Q(CACHE_ADDR2[1]) );
    zivb U1142 ( .A(CACHE_ADDR2[1]), .Y(n2183) );
    zdffqrb CACHE_ADDR2_reg_0 ( .CK(PCICLK), .D(CACHE_ADDR21034_0), .R(TRST_), 
        .Q(CACHE_ADDR2[0]) );
    zivb U1143 ( .A(CACHE_ADDR2[0]), .Y(n2181) );
    zdffqsb FROZEN_reg ( .CK(PCICLK), .D(FROZEN1654), .S(TRST_), .Q(FROZEN) );
    zdffqrb PERIODSM_reg_3 ( .CK(PCICLK), .D(PHASENXT_FetchTD), .R(TRST_), .Q(
        PERIODSM_3) );
    zivb U1144 ( .A(PERIODSM_3), .Y(n2229) );
    zdffrb EXEITD2_reg ( .CK(PCICLK), .D(EXEITD21109), .R(TRST_), .Q(EXEITD2), 
        .QN(n2409) );
    zdffqrb PERIODSM_reg_4 ( .CK(PCICLK), .D(PHASENXT_ParseTD), .R(TRST_), .Q(
        PHASE_ParseTD) );
    zivb U1145 ( .A(PHASE_ParseTD), .Y(n2228) );
    zdffqrb RECOVERYMODE_reg ( .CK(PCICLK), .D(RECOVERYMODE642), .R(TRST_), 
        .Q(RECOVERYMODE) );
    zivb U1146 ( .A(RECOVERYMODE), .Y(n2249) );
    zdffqrb TD_PARSE_GO2_T_reg ( .CK(PCICLK), .D(n2011), .R(TRST_), .Q(
        TD_PARSE_GO2_T) );
    zdffrb EXEQH2_reg ( .CK(PCICLK), .D(EXEQH21183), .R(TRST_), .Q(EXEQH2), 
        .QN(n2405) );
    zdffqrb DWNUM_reg_2 ( .CK(PCICLK), .D(DWNUM1434_2), .R(TRST_), .Q(DWNUM[2]
        ) );
    zdffqrb DWNUM_reg_3 ( .CK(PCICLK), .D(DWNUM1434_3), .R(TRST_), .Q(DWNUM[3]
        ) );
    zdffrb EXESITD1_reg ( .CK(PCICLK), .D(EXESITD11220), .R(TRST_), .Q(
        EXESITD1), .QN(n2403) );
    zdffqrb PERIODSM_reg_5 ( .CK(PCICLK), .D(PERIODSMNXT_5), .R(TRST_), .Q(
        PERIODSM_5) );
    zivb U1147 ( .A(PERIODSM_5), .Y(n2318) );
    zdffqrb PERIODSM_reg_2 ( .CK(PCICLK), .D(n2009), .R(TRST_), .Q(
        PHASE_FetchFSTN) );
    zivb U1148 ( .A(PHASE_FetchFSTN), .Y(n2245) );
    zdffqrb TRANEXED_reg ( .CK(PCICLK), .D(TRANEXED1556), .R(TRST_), .Q(
        TRANEXED) );
    zdffqrb TD_PARSE_GO1_T_reg ( .CK(PCICLK), .D(n2010), .R(TRST_), .Q(
        TD_PARSE_GO1_T) );
    zdffqrb CACHE_SEL_reg ( .CK(PCICLK), .D(CACHE_SEL_PRE), .R(TRST_), .Q(
        CACHE_SEL) );
    zivb U1149 ( .A(CACHE_SEL), .Y(n2023) );
    zdffrb EXEQH1_reg ( .CK(PCICLK), .D(EXEQH11146), .R(TRST_), .Q(EXEQH1), 
        .QN(n2407) );
    zdffrb PERIOD_RUN_reg ( .CK(PCICLK), .D(PERIOD_RUN_pre), .R(TRST_), .Q(
        PERIOD_RUN), .QN(n2140) );
    zdffrb EXEITD1_reg ( .CK(PCICLK), .D(EXEITD11072), .R(TRST_), .Q(EXEITD1), 
        .QN(n2411) );
    zdffqrb DWNUM_reg_1 ( .CK(PCICLK), .D(DWNUM1434_1), .R(TRST_), .Q(DWNUM[1]
        ) );
    zdffqsb EXE_HALT_reg ( .CK(PCICLK), .D(EXE_HALT_pre), .S(TRST_), .Q(
        EXE_HALT) );
    zdffrb EXESITD2_reg ( .CK(PCICLK), .D(EXESITD21257), .R(TRST_), .Q(
        EXESITD2), .QN(n2401) );
    zdffrb TD_ACT_SEL_reg ( .CK(PCICLK), .D(TD_ACT_SEL827), .R(TRST_), .Q(
        TD_ACT2), .QN(TD_ACT1) );
    zdffqsb DWNUM_reg_0 ( .CK(PCICLK), .D(DWNUM1434_0), .S(TRST_), .Q(DWNUM[0]
        ) );
    zdffrb PERIODSM_reg_6 ( .CK(PCICLK), .D(PERIODSMNXT_6), .R(TRST_), .Q(
        PERIODSM_6), .QN(n2172) );
    zdffqrb FRNUM_INC_reg ( .CK(PCICLK), .D(FRNUM_INC506), .R(TRST_), .Q(
        FRNUM_INC) );
    zivb U1150 ( .A(FRNUM_INC), .Y(n2357) );
    zdffqrb PERIODSM_reg_1 ( .CK(PCICLK), .D(PHASENXT_FetchPList), .R(TRST_), 
        .Q(PERIODSM_1) );
    zivb U1151 ( .A(PERIODSM_1), .Y(n2234) );
    zaoi21b U1152 ( .A(n2463), .B(n2464), .C(n2133), .Y(TDHCIGNT2) );
    zaoi21b U1153 ( .A(n2465), .B(n2466), .C(n2132), .Y(TDHCIGNT1) );
    znr2b U1154 ( .A(n2147), .B(n2231), .Y(n2009) );
    znr2b U1155 ( .A(PHASE_ParseTD), .B(n2241), .Y(n2010) );
    znr2b U1156 ( .A(PHASE_ParseTD), .B(n2240), .Y(n2011) );
    znr2b U1157 ( .A(LIST_SEL), .B(EHCIFLOW_IDLE), .Y(n2012) );
    znr4b U1158 ( .A(PERIOD_END), .B(PERIODSM_6), .C(n2228), .D(n2171), .Y(
        n2013) );
    znr3b U1159 ( .A(n2318), .B(n2168), .C(FETCHTD), .Y(n2014) );
    zaoi222b U1160 ( .A(n2348), .B(n2317), .C(n2122), .D(n2349), .E(TDIDLE1), 
        .F(n2160), .Y(n2015) );
    zivd U1161 ( .A(n2471), .Y(n2033) );
    zbfb U1162 ( .A(n2033), .Y(n2474) );
    zivb U1163 ( .A(n2361), .Y(n2016) );
    zivd U1164 ( .A(n2361), .Y(n2031) );
    zivb U1165 ( .A(n2368), .Y(n2017) );
    zivd U1166 ( .A(n2368), .Y(n2101) );
    zivb U1167 ( .A(n2364), .Y(n2018) );
    zao22b U1168 ( .A(n2030), .B(TDSTARTADR[7]), .C(n2016), .D(CACHE_ADDR2[2]), 
        .Y(CACHE_ADDR21034_2) );
    zao22b U1169 ( .A(n2030), .B(TDSTARTADR[11]), .C(n2031), .D(CACHE_ADDR2[6]
        ), .Y(CACHE_ADDR21034_6) );
    zao22b U1170 ( .A(n2030), .B(TDSTARTADR[18]), .C(n2016), .D(CACHE_ADDR2
        [13]), .Y(CACHE_ADDR21034_13) );
    zao22b U1171 ( .A(n2030), .B(TDSTARTADR[9]), .C(n2031), .D(CACHE_ADDR2[4]), 
        .Y(CACHE_ADDR21034_4) );
    zao22b U1172 ( .A(n2018), .B(TDSTARTADR[20]), .C(n2031), .D(CACHE_ADDR2
        [15]), .Y(CACHE_ADDR21034_15) );
    zao22b U1173 ( .A(n2030), .B(TDSTARTADR[22]), .C(n2031), .D(CACHE_ADDR2
        [17]), .Y(CACHE_ADDR21034_17) );
    zao22b U1174 ( .A(n2030), .B(TDSTARTADR[31]), .C(n2031), .D(CACHE_ADDR2
        [26]), .Y(CACHE_ADDR21034_26) );
    zao22b U1175 ( .A(n2030), .B(TDSTARTADR[13]), .C(n2031), .D(CACHE_ADDR2[8]
        ), .Y(CACHE_ADDR21034_8) );
    zao22b U1176 ( .A(n2018), .B(TDSTARTADR[30]), .C(n2031), .D(CACHE_ADDR2
        [25]), .Y(CACHE_ADDR21034_25) );
    zao22b U1177 ( .A(n2030), .B(TDSTARTADR[8]), .C(n2031), .D(CACHE_ADDR2[3]), 
        .Y(CACHE_ADDR21034_3) );
    zao22b U1178 ( .A(n2030), .B(TDSTARTADR[29]), .C(n2031), .D(CACHE_ADDR2
        [24]), .Y(CACHE_ADDR21034_24) );
    zao22b U1179 ( .A(n2030), .B(TDSTARTADR[24]), .C(n2031), .D(CACHE_ADDR2
        [19]), .Y(CACHE_ADDR21034_19) );
    zao22b U1180 ( .A(n2030), .B(TDSTARTADR[28]), .C(n2016), .D(CACHE_ADDR2
        [23]), .Y(CACHE_ADDR21034_23) );
    zao22b U1181 ( .A(n2030), .B(TDSTARTADR[14]), .C(n2031), .D(CACHE_ADDR2[9]
        ), .Y(CACHE_ADDR21034_9) );
    zao22b U1182 ( .A(n2030), .B(TDSTARTADR[27]), .C(n2016), .D(CACHE_ADDR2
        [22]), .Y(CACHE_ADDR21034_22) );
    zao22b U1183 ( .A(n2030), .B(TDSTARTADR[12]), .C(n2031), .D(CACHE_ADDR2[7]
        ), .Y(CACHE_ADDR21034_7) );
    zao22b U1184 ( .A(n2018), .B(TDSTARTADR[26]), .C(n2031), .D(CACHE_ADDR2
        [21]), .Y(CACHE_ADDR21034_21) );
    zao22b U1185 ( .A(n2030), .B(TDSTARTADR[10]), .C(n2031), .D(CACHE_ADDR2[5]
        ), .Y(CACHE_ADDR21034_5) );
    zao22b U1186 ( .A(n2030), .B(TDSTARTADR[25]), .C(n2016), .D(CACHE_ADDR2
        [20]), .Y(CACHE_ADDR21034_20) );
    zao22b U1187 ( .A(n2018), .B(TDSTARTADR[6]), .C(n2016), .D(CACHE_ADDR2[1]), 
        .Y(CACHE_ADDR21034_1) );
    zao22b U1188 ( .A(n2030), .B(TDSTARTADR[21]), .C(n2031), .D(CACHE_ADDR2
        [16]), .Y(CACHE_ADDR21034_16) );
    zao22b U1189 ( .A(n2018), .B(TDSTARTADR[23]), .C(n2016), .D(CACHE_ADDR2
        [18]), .Y(CACHE_ADDR21034_18) );
    zao22b U1190 ( .A(n2030), .B(TDSTARTADR[17]), .C(n2031), .D(CACHE_ADDR2
        [12]), .Y(CACHE_ADDR21034_12) );
    zao22b U1191 ( .A(n2018), .B(TDSTARTADR[19]), .C(n2031), .D(CACHE_ADDR2
        [14]), .Y(CACHE_ADDR21034_14) );
    zao22b U1192 ( .A(n2018), .B(TDSTARTADR[16]), .C(n2031), .D(CACHE_ADDR2
        [11]), .Y(CACHE_ADDR21034_11) );
    zao22b U1193 ( .A(n2018), .B(TDSTARTADR[5]), .C(n2016), .D(CACHE_ADDR2[0]), 
        .Y(CACHE_ADDR21034_0) );
    zao22b U1194 ( .A(n2030), .B(TDSTARTADR[15]), .C(n2031), .D(CACHE_ADDR2
        [10]), .Y(CACHE_ADDR21034_10) );
    zivd U1195 ( .A(n2364), .Y(n2030) );
    zivb U1196 ( .A(n2365), .Y(n2019) );
    zao22b U1197 ( .A(n2101), .B(TDSTARTADR[7]), .C(n2102), .D(CACHE_ADDR1[2]), 
        .Y(CACHE_ADDR1996_2) );
    zao22b U1198 ( .A(n2101), .B(TDSTARTADR[11]), .C(n2102), .D(CACHE_ADDR1[6]
        ), .Y(CACHE_ADDR1996_6) );
    zao22b U1199 ( .A(n2101), .B(TDSTARTADR[18]), .C(n2102), .D(CACHE_ADDR1
        [13]), .Y(CACHE_ADDR1996_13) );
    zao22b U1200 ( .A(n2101), .B(TDSTARTADR[9]), .C(n2102), .D(CACHE_ADDR1[4]), 
        .Y(CACHE_ADDR1996_4) );
    zao22b U1201 ( .A(n2017), .B(TDSTARTADR[20]), .C(n2019), .D(CACHE_ADDR1
        [15]), .Y(CACHE_ADDR1996_15) );
    zao22b U1202 ( .A(n2101), .B(TDSTARTADR[22]), .C(n2102), .D(CACHE_ADDR1
        [17]), .Y(CACHE_ADDR1996_17) );
    zao22b U1203 ( .A(n2101), .B(TDSTARTADR[31]), .C(n2102), .D(CACHE_ADDR1
        [26]), .Y(CACHE_ADDR1996_26) );
    zao22b U1204 ( .A(n2101), .B(TDSTARTADR[13]), .C(n2102), .D(CACHE_ADDR1[8]
        ), .Y(CACHE_ADDR1996_8) );
    zao22b U1205 ( .A(n2017), .B(TDSTARTADR[30]), .C(n2019), .D(CACHE_ADDR1
        [25]), .Y(CACHE_ADDR1996_25) );
    zao22b U1206 ( .A(n2101), .B(TDSTARTADR[8]), .C(n2102), .D(CACHE_ADDR1[3]), 
        .Y(CACHE_ADDR1996_3) );
    zao22b U1207 ( .A(n2101), .B(TDSTARTADR[29]), .C(n2102), .D(CACHE_ADDR1
        [24]), .Y(CACHE_ADDR1996_24) );
    zao22b U1208 ( .A(n2101), .B(TDSTARTADR[24]), .C(n2102), .D(CACHE_ADDR1
        [19]), .Y(CACHE_ADDR1996_19) );
    zao22b U1209 ( .A(n2101), .B(TDSTARTADR[28]), .C(n2102), .D(CACHE_ADDR1
        [23]), .Y(CACHE_ADDR1996_23) );
    zao22b U1210 ( .A(n2101), .B(TDSTARTADR[14]), .C(n2102), .D(CACHE_ADDR1[9]
        ), .Y(CACHE_ADDR1996_9) );
    zao22b U1211 ( .A(n2101), .B(TDSTARTADR[27]), .C(n2102), .D(CACHE_ADDR1
        [22]), .Y(CACHE_ADDR1996_22) );
    zao22b U1212 ( .A(n2101), .B(TDSTARTADR[12]), .C(n2102), .D(CACHE_ADDR1[7]
        ), .Y(CACHE_ADDR1996_7) );
    zao22b U1213 ( .A(n2017), .B(TDSTARTADR[26]), .C(n2019), .D(CACHE_ADDR1
        [21]), .Y(CACHE_ADDR1996_21) );
    zao22b U1214 ( .A(n2101), .B(TDSTARTADR[10]), .C(n2102), .D(CACHE_ADDR1[5]
        ), .Y(CACHE_ADDR1996_5) );
    zao22b U1215 ( .A(n2101), .B(TDSTARTADR[25]), .C(n2102), .D(CACHE_ADDR1
        [20]), .Y(CACHE_ADDR1996_20) );
    zao22b U1216 ( .A(n2017), .B(TDSTARTADR[6]), .C(n2019), .D(CACHE_ADDR1[1]), 
        .Y(CACHE_ADDR1996_1) );
    zao22b U1217 ( .A(n2101), .B(TDSTARTADR[21]), .C(n2102), .D(CACHE_ADDR1
        [16]), .Y(CACHE_ADDR1996_16) );
    zao22b U1218 ( .A(n2017), .B(TDSTARTADR[23]), .C(n2019), .D(CACHE_ADDR1
        [18]), .Y(CACHE_ADDR1996_18) );
    zao22b U1219 ( .A(n2101), .B(TDSTARTADR[17]), .C(n2102), .D(CACHE_ADDR1
        [12]), .Y(CACHE_ADDR1996_12) );
    zao22b U1220 ( .A(n2017), .B(TDSTARTADR[19]), .C(n2019), .D(CACHE_ADDR1
        [14]), .Y(CACHE_ADDR1996_14) );
    zao22b U1221 ( .A(n2017), .B(TDSTARTADR[16]), .C(n2019), .D(CACHE_ADDR1
        [11]), .Y(CACHE_ADDR1996_11) );
    zao22b U1222 ( .A(n2017), .B(TDSTARTADR[5]), .C(n2019), .D(CACHE_ADDR1[0]), 
        .Y(CACHE_ADDR1996_0) );
    zao22b U1223 ( .A(n2101), .B(TDSTARTADR[15]), .C(n2102), .D(CACHE_ADDR1
        [10]), .Y(CACHE_ADDR1996_10) );
    zivd U1224 ( .A(n2365), .Y(n2102) );
    zivb U1225 ( .A(n2027), .Y(n2020) );
    zoa211b U1226 ( .A(PHCI_DW0[0]), .B(n2155), .C(PCIEND), .D(n2156), .Y(
        n2110) );
    zor2b U1227 ( .A(n2112), .B(PCIEND), .Y(n2026) );
    zao32b U1228 ( .A(n2013), .B(n2129), .C(n2128), .D(PCIEND), .E(n2446), .Y(
        n2239) );
    zoa211b U1229 ( .A(PCIEND), .B(n2148), .C(n2149), .D(n2150), .Y(n2147) );
    zcxi5d U1230 ( .A(n2155), .B(n2316), .C(n2447), .D(PCIEND), .E(n2230), .Y(
        n2359) );
    zoa22b U1231 ( .A(n2104), .B(n2143), .C(n2020), .D(n2144), .Y(n2142) );
    zivb U1232 ( .A(PCIEND), .Y(n2027) );
    zdffsd PERIODSM_reg_0 ( .CK(PCICLK), .D(PERIODSMNXT_0), .S(TRST_), .Q(
        PERIOD_END), .QN(PERIOD_ACT) );
    zor3b U1233 ( .A(n2009), .B(PHASENXT_FetchTD), .C(PHASENXT_FetchPList), 
        .Y(FETCHTDNXT) );
    zan4b U1234 ( .A(TDIDLE2), .B(n2025), .C(TDIDLE1), .D(n2026), .Y(
        EXE_HALT_pre) );
    zao211b U1235 ( .A(FETCHTD), .B(n2027), .C(TDHCIGNT1), .D(TDHCIGNT2), .Y(
        EHCIREQ) );
    zao211b U1236 ( .A(TDSTARTADR[0]), .B(n2477), .C(n2037), .D(n2038), .Y(
        TDSTARTADR717_0) );
    zao211b U1237 ( .A(n2103), .B(n2104), .C(n2105), .D(n2106), .Y(
        PERIODSMNXT_0) );
    zoa21d U1238 ( .A(n2107), .B(n2108), .C(n2109), .Y(PERIODSMNXT_5) );
    zoa21d U1239 ( .A(n2110), .B(n2111), .C(n2109), .Y(PERIODSMNXT_6) );
    zao211b U1240 ( .A(DWNUM[0]), .B(n2112), .C(n2113), .D(n2009), .Y(
        DWNUM1434_0) );
    zao222b U1241 ( .A(FRNUM[12]), .B(n2117), .C(n2118), .D(FRNUM_PER_PRE_12), 
        .E(FRNUM_PER_PRE574_12), .F(n2119), .Y(FRNUM_PER_PRE597_12) );
    zao222b U1242 ( .A(FRNUM[11]), .B(n2117), .C(n2118), .D(FRNUM_PER_PRE_11), 
        .E(FRNUM_PER_PRE574_11), .F(n2119), .Y(FRNUM_PER_PRE597_11) );
    zao222b U1243 ( .A(n2118), .B(FRNUM_PER[10]), .C(FRNUM[10]), .D(n2117), 
        .E(FRNUM_PER_PRE574_10), .F(n2119), .Y(FRNUM_PER_PRE597_10) );
    zao222b U1244 ( .A(n2118), .B(FRNUM_PER[9]), .C(FRNUM[9]), .D(n2117), .E(
        n2119), .F(FRNUM_PER_PRE574_9), .Y(FRNUM_PER_PRE597_9) );
    zao222b U1245 ( .A(n2118), .B(FRNUM_PER[8]), .C(FRNUM[8]), .D(n2117), .E(
        FRNUM_PER_PRE574_8), .F(n2119), .Y(FRNUM_PER_PRE597_8) );
    zao222b U1246 ( .A(n2118), .B(FRNUM_PER[7]), .C(FRNUM[7]), .D(n2117), .E(
        FRNUM_PER_PRE574_7), .F(n2119), .Y(FRNUM_PER_PRE597_7) );
    zao222b U1247 ( .A(n2118), .B(FRNUM_PER[6]), .C(FRNUM[6]), .D(n2117), .E(
        FRNUM_PER_PRE574_6), .F(n2119), .Y(FRNUM_PER_PRE597_6) );
    zao222b U1248 ( .A(n2118), .B(FRNUM_PER[5]), .C(FRNUM[5]), .D(n2117), .E(
        FRNUM_PER_PRE574_5), .F(n2119), .Y(FRNUM_PER_PRE597_5) );
    zao222b U1249 ( .A(n2118), .B(FRNUM_PER[4]), .C(FRNUM[4]), .D(n2117), .E(
        FRNUM_PER_PRE574_4), .F(n2119), .Y(FRNUM_PER_PRE597_4) );
    zao222b U1250 ( .A(n2118), .B(FRNUM_PER[3]), .C(FRNUM[3]), .D(n2117), .E(
        FRNUM_PER_PRE574_3), .F(n2119), .Y(FRNUM_PER_PRE597_3) );
    zao222b U1251 ( .A(n2118), .B(FRNUM_PER[2]), .C(FRNUM[2]), .D(n2117), .E(
        FRNUM_PER_PRE574_2), .F(n2119), .Y(FRNUM_PER_PRE597_2) );
    zao222b U1252 ( .A(n2118), .B(FRNUM_PER[1]), .C(FRNUM[1]), .D(n2117), .E(
        FRNUM_PER_PRE574_1), .F(n2119), .Y(FRNUM_PER_PRE597_1) );
    zao222b U1253 ( .A(n2118), .B(FRNUM_PER[0]), .C(FRNUM[0]), .D(n2117), .E(
        FRNUM_PER_PRE574_0), .F(n2119), .Y(FRNUM_PER_PRE597_0) );
    zan4b U1254 ( .A(n2121), .B(n2114), .C(n2122), .D(n2123), .Y(n2120) );
    zan4b U1255 ( .A(RECOVERYMODE), .B(PERIOD_ACT), .C(n2134), .D(n2135), .Y(
        n2032) );
    zoa21d U1256 ( .A(n2152), .B(CACHEHIT1), .C(TDIDLE1), .Y(n2151) );
    zoa21d U1257 ( .A(n2152), .B(CACHEHIT2), .C(TDIDLE2), .Y(n2153) );
    zoa21d U1258 ( .A(n2154), .B(n2014), .C(n2157), .Y(n2111) );
    zoa21d U1259 ( .A(n2158), .B(n2014), .C(n2159), .Y(n2107) );
    zoa21d U1260 ( .A(PARSETDEND1), .B(PARSETDEND2), .C(n2013), .Y(n2108) );
    zoa21d U1261 ( .A(TDSTARTADR[1]), .B(n2116), .C(PHASENXT_FetchTD), .Y(
        n2113) );
    zor3b U1262 ( .A(n2196), .B(n2197), .C(n2198), .Y(n2199) );
    zor3b U1263 ( .A(n2193), .B(n2194), .C(n2195), .Y(n2200) );
    zor6b U1264 ( .A(n2201), .B(n2202), .C(n2203), .D(n2204), .E(n2205), .F(
        n2206), .Y(n2164) );
    zor6b U1265 ( .A(n2220), .B(n2221), .C(n2222), .D(n2223), .E(n2224), .F(
        n2225), .Y(n2162) );
    zor3b U1266 ( .A(n2170), .B(n2172), .C(n2171), .Y(n2227) );
    zor4b U1267 ( .A(n2229), .B(PERIODSM_5), .C(PCACHE_EN), .D(n2168), .Y(
        n2230) );
    zor3b U1268 ( .A(PERIODSM_3), .B(PERIODSM_5), .C(n2168), .Y(n2233) );
    zor3b U1269 ( .A(PHASE_FetchFSTN), .B(n2234), .C(n2233), .Y(n2144) );
    zor4b U1270 ( .A(PERIODSM_1), .B(PERIOD_END), .C(n2245), .D(n2027), .Y(
        n2246) );
    zor3b U1271 ( .A(n2244), .B(RECOVERYMODE), .C(PHCI_DW1[0]), .Y(n2247) );
    zor4b U1272 ( .A(n2249), .B(n2244), .C(n2250), .D(n2246), .Y(n2251) );
    zor4b U1273 ( .A(PERIOD_END), .B(PARSETDEND1), .C(n2129), .D(n2255), .Y(
        n2254) );
    zor3b U1274 ( .A(PERIOD_END), .B(n2128), .C(n2255), .Y(n2256) );
    zor4b U1275 ( .A(n2200), .B(n2339), .C(n2139), .D(n2199), .Y(n2104) );
    zor4b U1276 ( .A(PHASE_ParseTD), .B(PERIODSM_6), .C(PERIOD_ACT), .D(n2171), 
        .Y(n2143) );
    zor3b U1277 ( .A(PERIODSM_1), .B(n2245), .C(n2233), .Y(n2148) );
    zor3b U1278 ( .A(FRNUM_INC), .B(n2351), .C(n2339), .Y(n2352) );
    zor2d U1279 ( .A(n2353), .B(n2012), .Y(n2117) );
    zor3b U1280 ( .A(PERIOD_END), .B(CACHE_INVALID2), .C(n2362), .Y(n2361) );
    zor4b U1281 ( .A(TDSTARTADR[0]), .B(n2023), .C(n2348), .D(n2129), .Y(n2363
        ) );
    zor3b U1282 ( .A(PERIOD_END), .B(CACHE_INVALID2), .C(n2363), .Y(n2364) );
    zor3b U1283 ( .A(PERIOD_END), .B(CACHE_INVALID1), .C(n2366), .Y(n2365) );
    zor4b U1284 ( .A(TDSTARTADR[0]), .B(CACHE_SEL), .C(n2348), .D(n2128), .Y(
        n2367) );
    zor3b U1285 ( .A(PERIOD_END), .B(CACHE_INVALID1), .C(n2367), .Y(n2368) );
    zan4b U1286 ( .A(n2415), .B(n2416), .C(n2417), .D(n2317), .Y(n2414) );
    zan4b U1287 ( .A(n2419), .B(n2420), .C(n2421), .D(n2422), .Y(n2418) );
    zor4b U1288 ( .A(n2371), .B(n2372), .C(n2369), .D(n2370), .Y(n2429) );
    zor4b U1289 ( .A(n2373), .B(n2374), .C(n2375), .D(n2429), .Y(n2205) );
    zor4b U1290 ( .A(n2378), .B(n2379), .C(n2376), .D(n2377), .Y(n2204) );
    zan4b U1291 ( .A(n2431), .B(n2432), .C(n2433), .D(n2317), .Y(n2430) );
    zan4b U1292 ( .A(n2435), .B(n2436), .C(n2437), .D(n2438), .Y(n2434) );
    zor4b U1293 ( .A(n2382), .B(n2383), .C(n2380), .D(n2381), .Y(n2445) );
    zor4b U1294 ( .A(n2384), .B(n2385), .C(n2386), .D(n2445), .Y(n2224) );
    zor4b U1295 ( .A(n2389), .B(n2390), .C(n2387), .D(n2388), .Y(n2223) );
    zao222b U1296 ( .A(SAVEPTR_9), .B(n2448), .C(PHCI_DW1[9]), .D(n2449), .E(
        PHCI_DW0[9]), .F(n2482), .Y(n2055) );
    zao222b U1297 ( .A(n2131), .B(DW1_0[9]), .C(n2451), .D(DW2_0[9]), .E(
        TDSTARTADR[9]), .F(n2036), .Y(n2056) );
    zao222b U1298 ( .A(SAVEPTR_8), .B(n2480), .C(PHCI_DW1[8]), .D(n2483), .E(
        PHCI_DW0[8]), .F(n2450), .Y(n2053) );
    zao222b U1299 ( .A(DW1_0[8]), .B(n2131), .C(DW2_0[8]), .D(n2479), .E(
        TDSTARTADR[8]), .F(n2476), .Y(n2054) );
    zao222b U1300 ( .A(SAVEPTR_7), .B(n2448), .C(PHCI_DW1[7]), .D(n2449), .E(
        PHCI_DW0[7]), .F(n2481), .Y(n2051) );
    zao222b U1301 ( .A(DW1_0[7]), .B(n2478), .C(DW2_0[7]), .D(n2451), .E(
        TDSTARTADR[7]), .F(n2477), .Y(n2052) );
    zao222b U1302 ( .A(SAVEPTR_6), .B(n2480), .C(PHCI_DW1[6]), .D(n2483), .E(
        PHCI_DW0[6]), .F(n2482), .Y(n2049) );
    zao222b U1303 ( .A(DW1_0[6]), .B(n2131), .C(DW2_0[6]), .D(n2479), .E(
        TDSTARTADR[6]), .F(n2036), .Y(n2050) );
    zao222b U1304 ( .A(SAVEPTR_5), .B(n2448), .C(PHCI_DW1[5]), .D(n2449), .E(
        PHCI_DW0[5]), .F(n2450), .Y(n2047) );
    zao222b U1305 ( .A(DW1_0[5]), .B(n2478), .C(DW2_0[5]), .D(n2451), .E(
        TDSTARTADR[5]), .F(n2476), .Y(n2048) );
    zao222b U1306 ( .A(SAVEPTR_4), .B(n2480), .C(PHCI_DW1[4]), .D(n2483), .E(
        PHCI_DW0[4]), .F(n2481), .Y(n2045) );
    zao222b U1307 ( .A(DW2_0[4]), .B(n2479), .C(DW1_0[4]), .D(n2478), .E(
        TDSTARTADR[4]), .F(n2477), .Y(n2046) );
    zao222b U1308 ( .A(SAVEPTR_31), .B(n2448), .C(PHCI_DW1[31]), .D(n2449), 
        .E(PHCI_DW0[31]), .F(n2482), .Y(n2099) );
    zao222b U1309 ( .A(DW1_0[31]), .B(n2131), .C(DW2_0[31]), .D(n2479), .E(
        TDSTARTADR[31]), .F(n2036), .Y(n2100) );
    zao222b U1310 ( .A(SAVEPTR_30), .B(n2448), .C(PHCI_DW1[30]), .D(n2483), 
        .E(PHCI_DW0[30]), .F(n2450), .Y(n2097) );
    zao222b U1311 ( .A(DW1_0[30]), .B(n2478), .C(DW2_0[30]), .D(n2451), .E(
        TDSTARTADR[30]), .F(n2476), .Y(n2098) );
    zao222b U1312 ( .A(SAVEPTR_3), .B(n2480), .C(PHCI_DW1[3]), .D(n2449), .E(
        PHCI_DW0[3]), .F(n2481), .Y(n2043) );
    zao222b U1313 ( .A(DW2_0[3]), .B(n2451), .C(DW1_0[3]), .D(n2131), .E(
        TDSTARTADR[3]), .F(n2477), .Y(n2044) );
    zao222b U1314 ( .A(SAVEPTR_29), .B(n2480), .C(PHCI_DW1[29]), .D(n2483), 
        .E(PHCI_DW0[29]), .F(n2482), .Y(n2095) );
    zao222b U1315 ( .A(DW1_0[29]), .B(n2131), .C(DW2_0[29]), .D(n2479), .E(
        TDSTARTADR[29]), .F(n2036), .Y(n2096) );
    zao222b U1316 ( .A(SAVEPTR_28), .B(n2448), .C(PHCI_DW1[28]), .D(n2449), 
        .E(PHCI_DW0[28]), .F(n2450), .Y(n2093) );
    zao222b U1317 ( .A(DW1_0[28]), .B(n2478), .C(DW2_0[28]), .D(n2451), .E(
        TDSTARTADR[28]), .F(n2476), .Y(n2094) );
    zao222b U1318 ( .A(SAVEPTR_27), .B(n2448), .C(PHCI_DW1[27]), .D(n2483), 
        .E(PHCI_DW0[27]), .F(n2481), .Y(n2091) );
    zao222b U1319 ( .A(DW1_0[27]), .B(n2131), .C(DW2_0[27]), .D(n2479), .E(
        TDSTARTADR[27]), .F(n2477), .Y(n2092) );
    zao222b U1320 ( .A(SAVEPTR_26), .B(n2480), .C(PHCI_DW1[26]), .D(n2449), 
        .E(PHCI_DW0[26]), .F(n2482), .Y(n2089) );
    zao222b U1321 ( .A(DW1_0[26]), .B(n2478), .C(DW2_0[26]), .D(n2451), .E(
        TDSTARTADR[26]), .F(n2036), .Y(n2090) );
    zao222b U1322 ( .A(SAVEPTR_25), .B(n2480), .C(PHCI_DW1[25]), .D(n2483), 
        .E(PHCI_DW0[25]), .F(n2450), .Y(n2087) );
    zao222b U1323 ( .A(DW1_0[25]), .B(n2131), .C(DW2_0[25]), .D(n2479), .E(
        TDSTARTADR[25]), .F(n2476), .Y(n2088) );
    zao222b U1324 ( .A(SAVEPTR_24), .B(n2448), .C(PHCI_DW1[24]), .D(n2449), 
        .E(PHCI_DW0[24]), .F(n2481), .Y(n2085) );
    zao222b U1325 ( .A(DW1_0[24]), .B(n2478), .C(DW2_0[24]), .D(n2451), .E(
        TDSTARTADR[24]), .F(n2477), .Y(n2086) );
    zao222b U1326 ( .A(SAVEPTR_23), .B(n2480), .C(PHCI_DW1[23]), .D(n2483), 
        .E(PHCI_DW0[23]), .F(n2482), .Y(n2083) );
    zao222b U1327 ( .A(DW1_0[23]), .B(n2131), .C(DW2_0[23]), .D(n2479), .E(
        TDSTARTADR[23]), .F(n2036), .Y(n2084) );
    zao222b U1328 ( .A(SAVEPTR_22), .B(n2448), .C(PHCI_DW1[22]), .D(n2449), 
        .E(PHCI_DW0[22]), .F(n2450), .Y(n2081) );
    zao222b U1329 ( .A(DW1_0[22]), .B(n2478), .C(DW2_0[22]), .D(n2451), .E(
        TDSTARTADR[22]), .F(n2476), .Y(n2082) );
    zao222b U1330 ( .A(SAVEPTR_21), .B(n2480), .C(PHCI_DW1[21]), .D(n2483), 
        .E(PHCI_DW0[21]), .F(n2481), .Y(n2079) );
    zao222b U1331 ( .A(DW1_0[21]), .B(n2131), .C(DW2_0[21]), .D(n2479), .E(
        TDSTARTADR[21]), .F(n2477), .Y(n2080) );
    zao222b U1332 ( .A(SAVEPTR_20), .B(n2448), .C(PHCI_DW1[20]), .D(n2449), 
        .E(PHCI_DW0[20]), .F(n2482), .Y(n2077) );
    zao222b U1333 ( .A(DW1_0[20]), .B(n2478), .C(DW2_0[20]), .D(n2451), .E(
        TDSTARTADR[20]), .F(n2036), .Y(n2078) );
    zao222b U1334 ( .A(SAVEPTR_2), .B(n2480), .C(PHCI_DW1[2]), .D(n2483), .E(
        PHCI_DW0[2]), .F(n2450), .Y(n2041) );
    zao222b U1335 ( .A(DW1_0[2]), .B(n2131), .C(DW2_0[2]), .D(n2479), .E(
        TDSTARTADR[2]), .F(n2476), .Y(n2042) );
    zao222b U1336 ( .A(SAVEPTR_19), .B(n2448), .C(PHCI_DW1[19]), .D(n2449), 
        .E(PHCI_DW0[19]), .F(n2481), .Y(n2075) );
    zao222b U1337 ( .A(DW1_0[19]), .B(n2478), .C(DW2_0[19]), .D(n2451), .E(
        TDSTARTADR[19]), .F(n2477), .Y(n2076) );
    zao222b U1338 ( .A(SAVEPTR_18), .B(n2480), .C(PHCI_DW1[18]), .D(n2483), 
        .E(PHCI_DW0[18]), .F(n2482), .Y(n2073) );
    zao222b U1339 ( .A(DW1_0[18]), .B(n2131), .C(DW2_0[18]), .D(n2479), .E(
        TDSTARTADR[18]), .F(n2036), .Y(n2074) );
    zao222b U1340 ( .A(SAVEPTR_17), .B(n2448), .C(PHCI_DW1[17]), .D(n2449), 
        .E(PHCI_DW0[17]), .F(n2450), .Y(n2071) );
    zao222b U1341 ( .A(DW1_0[17]), .B(n2478), .C(DW2_0[17]), .D(n2451), .E(
        TDSTARTADR[17]), .F(n2476), .Y(n2072) );
    zao222b U1342 ( .A(SAVEPTR_16), .B(n2480), .C(PHCI_DW1[16]), .D(n2483), 
        .E(PHCI_DW0[16]), .F(n2481), .Y(n2069) );
    zao222b U1343 ( .A(DW1_0[16]), .B(n2131), .C(DW2_0[16]), .D(n2479), .E(
        TDSTARTADR[16]), .F(n2477), .Y(n2070) );
    zao222b U1344 ( .A(SAVEPTR_15), .B(n2448), .C(PHCI_DW1[15]), .D(n2449), 
        .E(PHCI_DW0[15]), .F(n2482), .Y(n2067) );
    zao222b U1345 ( .A(DW1_0[15]), .B(n2478), .C(DW2_0[15]), .D(n2451), .E(
        TDSTARTADR[15]), .F(n2036), .Y(n2068) );
    zao222b U1346 ( .A(SAVEPTR_14), .B(n2480), .C(PHCI_DW1[14]), .D(n2483), 
        .E(PHCI_DW0[14]), .F(n2450), .Y(n2065) );
    zao222b U1347 ( .A(DW1_0[14]), .B(n2131), .C(DW2_0[14]), .D(n2479), .E(
        TDSTARTADR[14]), .F(n2476), .Y(n2066) );
    zao222b U1348 ( .A(SAVEPTR_13), .B(n2448), .C(PHCI_DW1[13]), .D(n2449), 
        .E(PHCI_DW0[13]), .F(n2481), .Y(n2063) );
    zao222b U1349 ( .A(DW1_0[13]), .B(n2478), .C(DW2_0[13]), .D(n2451), .E(
        TDSTARTADR[13]), .F(n2477), .Y(n2064) );
    zao222b U1350 ( .A(SAVEPTR_12), .B(n2480), .C(PHCI_DW1[12]), .D(n2483), 
        .E(PHCI_DW0[12]), .F(n2482), .Y(n2061) );
    zao222b U1351 ( .A(DW1_0[12]), .B(n2131), .C(DW2_0[12]), .D(n2479), .E(
        TDSTARTADR[12]), .F(n2036), .Y(n2062) );
    zao222b U1352 ( .A(SAVEPTR_11), .B(n2448), .C(PHCI_DW1[11]), .D(n2449), 
        .E(PHCI_DW0[11]), .F(n2450), .Y(n2059) );
    zao222b U1353 ( .A(DW1_0[11]), .B(n2478), .C(DW2_0[11]), .D(n2451), .E(
        TDSTARTADR[11]), .F(n2476), .Y(n2060) );
    zao222b U1354 ( .A(SAVEPTR_10), .B(n2480), .C(PHCI_DW1[10]), .D(n2483), 
        .E(PHCI_DW0[10]), .F(n2481), .Y(n2057) );
    zao222b U1355 ( .A(DW1_0[10]), .B(n2131), .C(DW2_0[10]), .D(n2479), .E(
        TDSTARTADR[10]), .F(n2476), .Y(n2058) );
    zao222b U1356 ( .A(SAVEPTR_1), .B(n2448), .C(PHCI_DW1[1]), .D(n2449), .E(
        PHCI_DW0[1]), .F(n2482), .Y(n2039) );
    zao222b U1357 ( .A(DW1_0[1]), .B(n2478), .C(DW2_0[1]), .D(n2451), .E(
        TDSTARTADR[1]), .F(n2036), .Y(n2040) );
    zao222b U1358 ( .A(DW2_0[0]), .B(n2479), .C(SAVEPTR_0), .D(n2480), .E(
        PHCI_DW0[0]), .F(n2450), .Y(n2038) );
    zan4b U1359 ( .A(n2453), .B(n2454), .C(n2455), .D(n2456), .Y(n2452) );
    zan4b U1360 ( .A(n2457), .B(n2458), .C(n2459), .D(n2452), .Y(n2347) );
    zao222b U1361 ( .A(PHCI_DW0[0]), .B(n2447), .C(PERIODSM_6), .D(n2170), .E(
        PERIODSM_5), .F(FETCHTD), .Y(n2460) );
    zor4b U1362 ( .A(n2167), .B(n2461), .C(n2231), .D(n2460), .Y(n2106) );
    zao222b U1363 ( .A(PHASE_FetchFSTN), .B(PERIODSM_1), .C(PERIODSM_3), .D(
        PCACHE_EN), .E(PHASE_ParseTD), .F(PERIOD_END), .Y(n2461) );
    zind2d U1364 ( .A(n2339), .B(HCI_PRESOF), .Y(n2135) );
    zor5b U1365 ( .A(CACHE_HIT), .B(n2348), .C(n2227), .D(n2226), .E(n2393), 
        .Y(n2360) );
    zao211b U1366 ( .A(n2358), .B(n2238), .C(n2394), .D(n2172), .Y(n2166) );
    zor2d U1367 ( .A(n2127), .B(PERIOD_END), .Y(n2036) );
    zao32d U1368 ( .A(PERIODSM_1), .B(PERIOD_ACT), .C(PCIEND), .D(n2467), .E(
        n2469), .Y(n2450) );
    zor3b U1369 ( .A(PHASE_ParseTD), .B(n2318), .C(n2413), .Y(n2464) );
    zor3b U1370 ( .A(PHASE_ParseTD), .B(n2318), .C(n2470), .Y(n2466) );
    zor4b U1371 ( .A(n2245), .B(n2247), .C(PERIOD_END), .D(n2027), .Y(n2471)
         );
    zor4b U1372 ( .A(n2245), .B(n2244), .C(n2250), .D(n2027), .Y(n2134) );
    zor3b U1373 ( .A(FRNUM[0]), .B(FRNUM[1]), .C(FRNUM[2]), .Y(n2138) );
    zor4b U1374 ( .A(TDSTARTADR[0]), .B(n2114), .C(n2227), .D(n2145), .Y(n2150
        ) );
    zao211b U1375 ( .A(n2148), .B(n2237), .C(PHCI_DW0[0]), .D(n2155), .Y(n2149
        ) );
    zor3b U1376 ( .A(EXEQH2), .B(EXESITD2), .C(EXEITD2), .Y(n2021) );
    zor3b U1377 ( .A(EXEQH1), .B(EXESITD1), .C(EXEITD1), .Y(n2024) );
    zoai22d U1378 ( .A(n2339), .B(n2351), .C(n2012), .D(n2357), .Y(n2034) );
    zor3b U1379 ( .A(TDSTARTADR[1]), .B(n2116), .C(n2240), .Y(n2402) );
    zor3b U1380 ( .A(TDSTARTADR[1]), .B(n2116), .C(n2241), .Y(n2404) );
    zor3b U1381 ( .A(TDSTARTADR[2]), .B(n2115), .C(n2240), .Y(n2406) );
    zor3b U1382 ( .A(TDSTARTADR[2]), .B(n2115), .C(n2241), .Y(n2408) );
    zor3b U1383 ( .A(TDSTARTADR[1]), .B(TDSTARTADR[2]), .C(n2240), .Y(n2410)
         );
    zor3b U1384 ( .A(TDSTARTADR[1]), .B(TDSTARTADR[2]), .C(n2241), .Y(n2412)
         );
    zor2d U1385 ( .A(n2127), .B(PERIOD_END), .Y(n2476) );
    zor2d U1386 ( .A(n2127), .B(PERIOD_END), .Y(n2477) );
    zao32d U1387 ( .A(PERIODSM_1), .B(PERIOD_ACT), .C(PCIEND), .D(n2467), .E(
        n2469), .Y(n2481) );
    zao32d U1388 ( .A(PERIODSM_1), .B(PERIOD_ACT), .C(PCIEND), .D(n2467), .E(
        n2469), .Y(n2482) );
endmodule


module PQHCTL ( QH_PARSE_GO, PARSEQHEND, QHPARSING, QHIDLE, FRNUM, DW0, DW1, 
    DW2, DW3, DW4, DW5, DW6, DW7, DW8, DW9, DW10, DW11, GEN_PERR, PCIEND, 
    UP_DW3, UP_DW6, UP_DW7, UP_DW8, UP_DW9, UP_LDW3, UP_LDW6, UP_LDW7, UP_LDW8, 
    UP_LDW9, CACHEPHASE, QHCIREQ, QHDWNUM, QDWOFFSET, QHCIADR, QHCIADD, 
    QHCIMWR, DWCNT, QHSM, TRAN_CMD, QH_ACT, QBUI_GO, CACHE_ADDR, CACHE_INVALID, 
    CRCERR, ACTLEN, BABBLE, PIDERR, TMOUT, RXNAK, RXNYET, RXSTALL, RXACK, 
    RXDATA0, RXDATA1, RXMDATA, RXPIDERR, TOGMATCH, SPD, EHCI_MAC_EOT, FEMPTY, 
    TDMAEND, QRXERR, HCI_PRESOF, MAXLEN, QCMDSTART_REQ, QCMDSTART, QEOT, 
    QTDEXE, LTINT_PCLK, USBINT_EN, ERRINT_EN, USBINT, ERRINT, QHIOCINT_S, 
    QHERRINT_S, QHIOCINT, QHERRINT, RECOVERYMODE, PCICLK, EHCIFLOW_PCLK, TRST_
     );
input  [13:0] FRNUM;
input  [31:0] DW0;
input  [31:0] DW7;
input  [31:0] DW9;
output [31:0] UP_DW8;
output [31:0] UP_DW6;
output [3:0] QDWOFFSET;
input  [26:0] CACHE_ADDR;
input  [31:0] DW1;
input  [31:0] DW6;
output [31:0] UP_DW7;
output [31:0] UP_DW9;
output [13:0] QHSM;
input  [31:0] DW2;
input  [31:0] DW3;
input  [31:0] DW8;
input  [3:0] DWCNT;
input  [31:0] DW4;
output [31:0] QHCIADR;
output [31:0] QHCIADD;
input  [10:0] ACTLEN;
input  [31:0] DW5;
input  [31:0] DW10;
input  [31:0] DW11;
output [104:0] TRAN_CMD;
output [10:0] MAXLEN;
output [31:0] UP_DW3;
output [3:0] QHDWNUM;
input  QH_PARSE_GO, GEN_PERR, PCIEND, QH_ACT, CRCERR, BABBLE, PIDERR, TMOUT, 
    RXNAK, RXNYET, RXSTALL, RXACK, RXDATA0, RXDATA1, RXMDATA, RXPIDERR, 
    TOGMATCH, SPD, EHCI_MAC_EOT, FEMPTY, TDMAEND, HCI_PRESOF, QCMDSTART, 
    LTINT_PCLK, USBINT_EN, ERRINT_EN, USBINT, ERRINT, RECOVERYMODE, PCICLK, 
    EHCIFLOW_PCLK, TRST_;
output PARSEQHEND, QHPARSING, QHIDLE, UP_LDW3, UP_LDW6, UP_LDW7, UP_LDW8, 
    UP_LDW9, CACHEPHASE, QHCIREQ, QHCIMWR, QBUI_GO, CACHE_INVALID, QRXERR, 
    QCMDSTART_REQ, QEOT, QTDEXE, QHIOCINT_S, QHERRINT_S, QHIOCINT, QHERRINT;
    wire VIR_TOTALBYTES_9, TOTALBYTES792_5, PING_ERR1014, OVERWBOFFSET2136_1, 
        VIR_TOTALBYTES_13, OVERWBOFFSET_P2090_5, SBYTES966_5, CURQTDPTR1736_27, 
        SPAREO6, HCI_PRESOF_T, MULT_1, SBYTES962_3, MINUEND_8, CPAGE1173_1, 
        XACTERR1308, TOTALBYTES_12, TOTALBYTES_6, TOTALBYTES_REAL_5, QHSMNXT_8, 
        PARSEQHEND_PRE, FRAMETAG1498_3, VIR_TOTALBYTES_0, OVERWBOFFSET2136_8, 
        TOTAL_SBYTES_14, TOTALBYTES792_14, TOTAL_SBYTES_2, 
        OVERWBOFFSET_P2070_2, QHSMNXT_12, CURQTDPTR1736_7, MULT588_0, 
        CPROGMASK1402_3, CURQTDPTR1736_12, CPAGE_0, QCMDSTART_EOT2265, 
        QHSMNXT_1, TOTALBYTES_8, NXTISSTSWB, MINUEND_6, TOTALBYTES_REAL_11, 
        FRAMETAG1470_2, CURQTDPTR1736_15, SPAREO0_, CPROGMASK1402_4, 
        CURQTDPTR1736_29, OVERWBOFFSET_P2070_5, SPAREO8, VIR_TOTALBYTES_7, 
        TOTAL_SBYTES_5, TOTALBYTES792_13, MINUEND_10, TOTAL_SBYTES_13, 
        TOTALBYTES_1, FRAMETAG1498_4, TOTALBYTES_REAL_2, SBYTES962_4, 
        CURQTDPTR1736_20, SBYTES966_2, VIR_TOTALBYTES_14, QHERRINT_T2413, 
        CURQTDPTR1736_9, OVERWBOFFSET_P2090_2, SPAREO1, OVERWBOFFSET2136_6, 
        TOTALBYTES792_2, VIR_TOTALBYTES_6, TOTAL_SBYTES_4, TOTALBYTES792_12, 
        TOTAL_SBYTES_12, CURQTDPTR1736_28, OVERWBOFFSET_P2070_4, UP_CACHE1, 
        SPAREO9, QCMDSTART_EOT, PHASENXT_resultwb, MINUEND_7, FRAMETAG1470_3, 
        CURQTDPTR1736_14, PHASENXT_idle, CPROGMASK1402_5, IMMEDRETRY, 
        TOTALBYTES_9, QHSMNXT_7, CUROFFSET_T_12, LENGTMAX867, 
        OVERWBOFFSET2136_7, TOTALBYTES792_3, CURQTDPTR1736_21, CURQTDPTR1736_8, 
        OVERWBOFFSET_P2090_3, SBYTES966_3, QHIOCINT2376, CPAGE1177_1, SPAREO0, 
        SBYTES962_5, TOTALBYTES_0, CACHE_INVALID1964, TOTALBYTES_REAL_3, 
        TOTALBYTES_14, OVERWBOFFSET_P2070_12, CACHE_MODIFY502, TOTALBYTES_7, 
        TOTALBYTES_13, QHSMNXT_9, TOTALBYTES_REAL_4, FRAMETAG1498_2, 
        SBYTES962_2, MULT_0, QRXERR_CUR1646, MINUEND_9, CPAGE1173_0, 
        SBYTES966_4, VIR_TOTALBYTES_12, OVERWBOFFSET_P2090_4, CURQTDPTR1736_26, 
        SPAREO7, VIR_TOTALBYTES_8, QHSM_12, DT1086, TOTALBYTES792_4, 
        OVERWBOFFSET2136_0, CPAGE_1, OVERWBOFFSET_P2090_12, CPROGMASK1402_2, 
        CURQTDPTR1736_13, FRAMETAG1470_4, OVERWBOFFSET_P2070_3, QHSMNXT_13, 
        CURQTDPTR1736_6, MULT588_1, QHIOCINT_T2339, VIR_TOTALBYTES_1, 
        OVERWBOFFSET2136_9, TOTAL_SBYTES_3, OVERWBOFFSET2136_2, TOTAL_SBYTES_8, 
        INACT_COND, TOTALBYTES792_6, ACTIVE, ACTIVE_NXT, QTDHALT, 
        OVERWBOFFSET2136_10, DT, SPAREO5, OVERWBOFFSET_P2070_8, 
        VIR_TOTALBYTES_10, OVERWBOFFSET_P2090_6, SBYTES966_6, CURQTDPTR1736_24, 
        CPAGE1173_2, CURQTDPTR1736_18, SBYTES962_0, FRAMETAG1498_0, 
        TOTALBYTES_11, TOTALBYTES_REAL_6, TOTALBYTES_5, SPLITXSTATE_OLD1378, 
        OVERWBOFFSET_P2070_10, TOTAL_SBYTES_1, VIR_TOTALBYTES_3, 
        OVERWBOFFSET_P2070_1, CURQTDPTR1736_11, CPROGMASK1402_0, MULT572_1, 
        QHSMNXT_2, OVERWBOFFSET_P2090_10, QHSMNXT_5, TOTALBYTES_REAL_8, 
        CURQTDPTR1736_31, CERR1251_1, CPROGMASK1402_7, FRAMETAG1470_1, 
        CURQTDPTR1736_16, MINUEND_5, TOTALBYTES_REAL_12, QHIOCINT_T, 
        OVERWBOFFSET_P2070_6, SPLITXSTATE1341, OVERWBOFFSET_P2090_8, 
        ACCEPT_DATA, QHERRINT2450, TOTAL_SBYTES_10, IMMEDRETRY1571, 
        TOTAL_SBYTES_6, TOTALBYTES792_10, VIR_TOTALBYTES_4, TOTALBYTES792_8, 
        TOTALBYTES_2, CERR_1, SPAREO2, CURQTDPTR1736_23, SBYTES966_1, 
        OVERWBOFFSET_P2090_1, TOTALBYTES792_1, OVERWBOFFSET2136_5, 
        TOTAL_SBYTES_11, TOTALBYTES792_11, TOTAL_SBYTES_7, TOTALBYTES792_9, 
        VIR_TOTALBYTES_5, QEOT2302, OVERWBOFFSET_P2070_7, LENGTMAX_PRE, 
        OVERWBOFFSET_P2090_9, CURQTDPTR1736_30, CPROGMASK1402_6, CERR1251_0, 
        FRAMETAG1470_0, CURQTDPTR1736_17, TOTALBYTES_REAL_13, MINUEND_4, 
        PHASENXT_outcyc, QHSMNXT_4, TOTALBYTES_REAL_9, TOTALBYTES792_0, 
        OVERWBOFFSET2136_4, CPAGE1177_2, SPAREO3, CURQTDPTR1736_22, SPAREO1_, 
        OVERWBOFFSET_P2090_0, SBYTES966_0, HCI_PRESOF_T1608, CERR_0, 
        SBYTES962_6, CACHE_MODIFY, TOTALBYTES_3, FRAMETAG1498_1, TOTALBYTES_10, 
        TOTALBYTES_REAL_7, TOTALBYTES_4, OVERWBOFFSET_P2070_11, LDPARM, 
        MISUF1318, CURQTDPTR1736_19, SBYTES962_1, SPAREO4, 
        OVERWBOFFSET_P2070_9, VIR_TOTALBYTES_11, OVERWBOFFSET_P2090_7, 
        CURQTDPTR1736_25, OVERWBOFFSET2136_3, TOTAL_SBYTES_9, TOTALBYTES792_7, 
        QHERRINT_T, OVERWBOFFSET2136_11, QHSMNXT_3, OVERWBOFFSET_P2090_11, 
        PING_ERR, CPAGE_2, CURQTDPTR1736_10, CPROGMASK1402_1, MINUEND_3, 
        MULT572_0, TOTALBYTES_REAL_14, CERR1255_1, CURQTDPTR1736_5, 
        OVERWBOFFSET_P2070_0, QHSMNXT_10, TOTAL_SBYTES_0, VIR_TOTALBYTES_2, 
        n2519, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, 
        n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, 
        n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2908, 
        n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, 
        n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, 
        n2930, n2931, n2932, n3023, n3029, n3030, n3031, n3032, n3033, n3034, 
        n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, 
        n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, 
        n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, 
        n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, 
        n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, 
        add_922_carry_8, add_922_carry_1, add_922_carry_7, add_922_carry_6, 
        add_922_carry_9, add_922_carry_2, add_922_carry_11, add_922_carry_10, 
        add_922_carry_5, add_922_carry_4, add_922_carry_3, sub_451_carry_1, 
        sub_451_carry_8, sub_451_carry_14, sub_451_carry_13, sub_451_carry_12, 
        sub_451_carry_7, sub_451_carry_6, sub_451_carry_9, sub_451_carry_2, 
        sub_451_carry_11, sub_451_carry_10, sub_451_carry_5, sub_451_carry_4, 
        sub_451_carry_3, sub_457_carry_1, sub_457_B_not_10, sub_457_B_not_8, 
        sub_457_carry_8, sub_457_B_not_6, sub_457_carry_14, sub_457_carry_13, 
        sub_457_carry_12, sub_457_carry_7, sub_457_carry_6, sub_457_B_not_7, 
        sub_457_B_not_9, sub_457_carry_9, sub_457_carry_2, sub_457_B_not_5, 
        sub_457_carry_11, sub_457_carry_10, sub_457_carry_5, sub_457_carry_4, 
        sub_457_B_not_4, sub_457_carry_3, sub_457_B_not_3, add_508_carry_1, 
        add_508_carry_6, add_508_carry_2, add_508_carry_5, add_508_carry_4, 
        add_508_carry_3, n3085, r469_carry_2, r469_carry_4, r469_carry_3, 
        add_919_carry_8, add_919_carry_1, add_919_carry_12, add_919_carry_7, 
        add_919_carry_6, add_919_carry_9, add_919_carry_2, add_919_carry_11, 
        add_919_carry_10, add_919_carry_5, add_919_carry_4, add_919_carry_3, 
        r481_carry_8, r481_carry_1, r481_carry_7, r481_carry_6, r481_carry_9, 
        r481_carry_2, r481_carry_11, r481_carry_10, r481_carry_5, r481_carry_4, 
        r481_carry_3, r489_carry_2, n3086, n3087, n3088, n3089, n3090, n3091, 
        n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
        n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, 
        n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
        n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
        n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, 
        n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, 
        n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, 
        n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, 
        n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, 
        n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, 
        n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
        n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
        n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, 
        n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, 
        n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, 
        n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, 
        n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, 
        n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, 
        n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, 
        n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, 
        n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, 
        n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, 
        n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, 
        n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, 
        n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, 
        n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, 
        n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, 
        n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, 
        n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, 
        n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, 
        n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, 
        n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, 
        n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, 
        n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, 
        n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, 
        n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, 
        n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, 
        n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, 
        n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, 
        n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, 
        n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, 
        n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, 
        n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, 
        n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, 
        n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, 
        n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, 
        n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, 
        n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, 
        n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, 
        n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, 
        n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, 
        n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, 
        n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, 
        n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, 
        n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, 
        n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, 
        n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, 
        n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, 
        n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, 
        n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, 
        n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, 
        n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, 
        n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, 
        n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, 
        n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, 
        n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, 
        n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, 
        n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, 
        n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, 
        n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, 
        n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, 
        n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, 
        n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, 
        n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, 
        n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, 
        n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, 
        n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, 
        n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, 
        n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, 
        n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, 
        n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, 
        n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, 
        n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, 
        n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, 
        n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, 
        n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, 
        n3952, n3953, n3954, n3955, n3956;
    assign UP_DW3[4] = 1'b0;
    assign UP_DW3[3] = 1'b0;
    assign UP_DW3[2] = 1'b0;
    assign UP_DW3[1] = 1'b0;
    assign UP_DW3[0] = 1'b0;
    assign UP_DW8[11] = 1'b0;
    assign UP_DW8[10] = 1'b0;
    assign UP_DW8[9] = 1'b0;
    assign UP_DW8[8] = 1'b0;
    assign QDWOFFSET[3] = 1'b0;
    assign QDWOFFSET[2] = 1'b1;
    assign QDWOFFSET[1] = 1'b0;
    assign QDWOFFSET[0] = 1'b0;
    assign QHCIADR[1] = 1'b0;
    assign QHCIADR[0] = 1'b0;
    assign TRAN_CMD[51] = 1'b0;
    assign TRAN_CMD[12] = 1'b0;
    assign TRAN_CMD[11] = 1'b1;
    assign TRAN_CMD[10] = 1'b1;
    assign TRAN_CMD[5] = 1'b0;
    assign TRAN_CMD[2] = 1'b0;
    zoai21b SPARE845 ( .A(SPAREO1), .B(LDPARM), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE842 ( .A(SPAREO0), .B(n2920), .C(SPAREO1_), .D(NXTISSTSWB), 
        .Y(SPAREO2) );
    zaoi211b SPARE843 ( .A(SPAREO4), .B(PARSEQHEND_PRE), .C(SPAREO6), .D(1'b0), 
        .Y(SPAREO8) );
    zoai21b SPARE844 ( .A(SPAREO0), .B(SPAREO8), .C(ACCEPT_DATA), .Y(SPAREO9)
         );
    znr3b SPARE846 ( .A(SPAREO2), .B(n2923), .C(SPAREO0_), .Y(SPAREO4) );
    zdffrb SPARE841 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE848 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE840 ( .CK(PCICLK), .D(INACT_COND), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE849 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb SPARE847 ( .A(SPAREO4), .Y(SPAREO5) );
    znd2b U892 ( .A(n2879), .B(n3082), .Y(n3049) );
    zivb U893 ( .A(DW1[17]), .Y(n3082) );
    zivb U894 ( .A(DW1[18]), .Y(n3056) );
    znd2b U895 ( .A(n2880), .B(n3051), .Y(n3080) );
    zivb U896 ( .A(DW1[16]), .Y(n3051) );
    znd2b U897 ( .A(TOTALBYTES_REAL_3), .B(n3055), .Y(n3045) );
    zivb U898 ( .A(DW1[19]), .Y(n3055) );
    znd2b U899 ( .A(TOTALBYTES_REAL_4), .B(n3057), .Y(n3046) );
    zivb U900 ( .A(DW1[20]), .Y(n3057) );
    znd2b U901 ( .A(n3048), .B(n3047), .Y(n3076) );
    znd2b U902 ( .A(DW1[19]), .B(n3916), .Y(n3048) );
    znd2b U903 ( .A(DW1[18]), .B(n3917), .Y(n3047) );
    znr2b U904 ( .A(n3083), .B(n3080), .Y(n3081) );
    znd2b U905 ( .A(TOTALBYTES_REAL_5), .B(n3054), .Y(n3041) );
    zivb U906 ( .A(DW1[21]), .Y(n3054) );
    znd2b U907 ( .A(TOTALBYTES_REAL_6), .B(n3058), .Y(n3042) );
    zivb U908 ( .A(DW1[22]), .Y(n3058) );
    znd2b U909 ( .A(n3044), .B(n3043), .Y(n3072) );
    znd2b U910 ( .A(DW1[21]), .B(n3914), .Y(n3044) );
    znd2b U911 ( .A(DW1[20]), .B(n3915), .Y(n3043) );
    znd2b U912 ( .A(n3046), .B(n3045), .Y(n3074) );
    zan2b U913 ( .A(n3526), .B(n3527), .Y(n3525) );
    znd2b U914 ( .A(TOTALBYTES_REAL_7), .B(n3053), .Y(n3037) );
    zivb U915 ( .A(DW1[23]), .Y(n3053) );
    znd2b U916 ( .A(TOTALBYTES_REAL_8), .B(n3059), .Y(n3038) );
    zivb U917 ( .A(DW1[24]), .Y(n3059) );
    znd2b U918 ( .A(n3040), .B(n3039), .Y(n3068) );
    znd2b U919 ( .A(DW1[23]), .B(n3912), .Y(n3040) );
    znd2b U920 ( .A(DW1[22]), .B(n3913), .Y(n3039) );
    znr2b U921 ( .A(n3073), .B(n3070), .Y(n3071) );
    znr2b U922 ( .A(n3075), .B(n3072), .Y(n3073) );
    znd2b U923 ( .A(n3042), .B(n3041), .Y(n3070) );
    zxo2b U924 ( .A(n3502), .B(n3822), .Y(n3694) );
    zxo2b U925 ( .A(n3500), .B(n3821), .Y(n3695) );
    zxo2b U926 ( .A(n3506), .B(n3820), .Y(n3696) );
    zivb U927 ( .A(DW2[11]), .Y(n3506) );
    zxo2b U928 ( .A(n3510), .B(n3819), .Y(n3697) );
    zivb U929 ( .A(DW2[9]), .Y(n3510) );
    zxo2b U930 ( .A(DW2[8]), .B(n3525), .Y(n3698) );
    zoai2x4b U931 ( .A(n3662), .B(n3670), .C(n3659), .D(n3669), .E(n3527), .F(
        n3526), .G(n3603), .H(n3668), .Y(n3672) );
    zoai2x4b U932 ( .A(n3658), .B(n3664), .C(n3660), .D(n3665), .E(n3663), .F(
        n3667), .G(n3661), .H(n3666), .Y(n3671) );
    zxo2b U933 ( .A(UP_DW9[2]), .B(FRNUM[5]), .Y(n3677) );
    zxo2b U934 ( .A(UP_DW9[4]), .B(FRNUM[7]), .Y(n3676) );
    zxo2b U935 ( .A(FRNUM[3]), .B(UP_DW9[0]), .Y(n3675) );
    zxo2b U936 ( .A(UP_DW9[3]), .B(FRNUM[6]), .Y(n3674) );
    zxo2b U937 ( .A(UP_DW9[1]), .B(FRNUM[4]), .Y(n3673) );
    znd2b U938 ( .A(n2878), .B(n3060), .Y(n3033) );
    znd2b U939 ( .A(TOTALBYTES_REAL_9), .B(n3052), .Y(n3034) );
    zivb U940 ( .A(DW1[25]), .Y(n3052) );
    znd2b U941 ( .A(n3036), .B(n3035), .Y(n3064) );
    znd2b U942 ( .A(DW1[25]), .B(n3910), .Y(n3036) );
    znd2b U943 ( .A(DW1[24]), .B(n3911), .Y(n3035) );
    znr2b U944 ( .A(n3069), .B(n3066), .Y(n3067) );
    znr2b U945 ( .A(n3071), .B(n3068), .Y(n3069) );
    znd2b U946 ( .A(n3038), .B(n3037), .Y(n3066) );
    zoai2x4b U947 ( .A(n3660), .B(n3504), .C(n3659), .D(n3502), .E(n3658), .F(
        n3500), .G(n3603), .H(n3514), .Y(n3679) );
    zivb U948 ( .A(DW2[12]), .Y(n3504) );
    zivb U949 ( .A(DW2[13]), .Y(n3502) );
    zivb U950 ( .A(DW2[14]), .Y(n3500) );
    zivb U951 ( .A(DW2[15]), .Y(n3514) );
    zivc U952 ( .A(n3660), .Y(n3351) );
    zivc U953 ( .A(n3659), .Y(n3352) );
    zoai2x4b U954 ( .A(n3527), .B(n3688), .C(n3663), .D(n3687), .E(n3662), .F(
        n3686), .G(n3661), .H(n3685), .Y(n3846) );
    zivb U955 ( .A(DW2[0]), .Y(n3688) );
    zivb U956 ( .A(n3527), .Y(n3346) );
    zivc U957 ( .A(n3663), .Y(n3348) );
    zivc U958 ( .A(n3662), .Y(n3349) );
    zivc U959 ( .A(n3661), .Y(n3350) );
    zoai2x4b U960 ( .A(n3690), .B(n3775), .C(n3654), .D(n3595), .E(n3855), .F(
        n3856), .G(n3857), .H(n3858), .Y(n3854) );
    znd8b U961 ( .A(n3715), .B(n3721), .C(n3719), .D(n3726), .E(n3723), .F(
        n3728), .G(n3730), .H(n3732), .Y(n3568) );
    zivb U962 ( .A(RXACK), .Y(n3546) );
    zivb U963 ( .A(RXNYET), .Y(n3699) );
    znd8b U964 ( .A(n3760), .B(n3761), .C(n3759), .D(n3757), .E(n3758), .F(
        n3756), .G(n3763), .H(n3762), .Y(n3618) );
    zivb U965 ( .A(TOGMATCH), .Y(n3627) );
    zor2b U966 ( .A(n2875), .B(n2873), .Y(n3848) );
    znr6b U967 ( .A(RXPIDERR), .B(RXACK), .C(RXNYET), .D(RXSTALL), .E(RXNAK), 
        .F(TOGMATCH), .Y(n3494) );
    zor2b U968 ( .A(QHSM[9]), .B(QHSM[11]), .Y(n3573) );
    zivb U969 ( .A(n3645), .Y(n3857) );
    znr2b U970 ( .A(n2878), .B(n3060), .Y(n3061) );
    zivb U971 ( .A(DW1[26]), .Y(n3060) );
    znr2b U972 ( .A(n3065), .B(n3062), .Y(n3063) );
    znr2b U973 ( .A(n3067), .B(n3064), .Y(n3065) );
    znd2b U974 ( .A(n3034), .B(n3033), .Y(n3062) );
    znd2b U975 ( .A(n3031), .B(n3030), .Y(n3032) );
    zivb U976 ( .A(DW9[7]), .Y(n3539) );
    zivb U977 ( .A(DW9[11]), .Y(n3540) );
    zivb U978 ( .A(DW9[6]), .Y(n3541) );
    zivb U979 ( .A(DW9[9]), .Y(n3635) );
    zivb U980 ( .A(DW9[8]), .Y(n3636) );
    zivb U981 ( .A(DW9[10]), .Y(n3634) );
    zivb U982 ( .A(DW9[5]), .Y(n3637) );
    zan2b U983 ( .A(n3519), .B(n3560), .Y(n3559) );
    zivb U984 ( .A(n3678), .Y(n3519) );
    zor2b U985 ( .A(n3126), .B(n3523), .Y(n3563) );
    zan2b U986 ( .A(n3583), .B(n3584), .Y(n3582) );
    zor2b U987 ( .A(n3638), .B(n3645), .Y(n3646) );
    znd2b U988 ( .A(n3583), .B(n3924), .Y(n3836) );
    zivb U989 ( .A(n3646), .Y(n3584) );
    zor2b U990 ( .A(n3106), .B(n3532), .Y(n3638) );
    zivb U991 ( .A(n3638), .Y(n3858) );
    zivb U992 ( .A(n3651), .Y(n3583) );
    zmux21lb U993 ( .A(CERR_1), .B(CERR1255_1), .S(n3923), .Y(n3612) );
    zxo2b U994 ( .A(n3085), .B(CERR_0), .Y(CERR1255_1) );
    zmux21lb U995 ( .A(CERR_0), .B(n3828), .S(n3923), .Y(n3615) );
    zoa22b U996 ( .A(QHSM[6]), .B(n3113), .C(QHSM[8]), .D(n3112), .Y(n3598) );
    zan2b U997 ( .A(TOTAL_SBYTES_14), .B(n3329), .Y(TOTALBYTES_REAL_14) );
    zan2b U998 ( .A(TOTAL_SBYTES_13), .B(n3329), .Y(TOTALBYTES_REAL_13) );
    zan2b U999 ( .A(TOTAL_SBYTES_12), .B(n3329), .Y(TOTALBYTES_REAL_12) );
    zivb U1000 ( .A(TOTALBYTES_REAL_12), .Y(n3030) );
    zan2b U1001 ( .A(TOTAL_SBYTES_11), .B(n3329), .Y(TOTALBYTES_REAL_11) );
    zivb U1002 ( .A(TOTALBYTES_REAL_11), .Y(n3031) );
    zor2b U1003 ( .A(TRAN_CMD[14]), .B(n3658), .Y(n3604) );
    zivd U1004 ( .A(n3658), .Y(n3353) );
    zor2b U1005 ( .A(n3753), .B(n3631), .Y(n3767) );
    zor2b U1006 ( .A(n3567), .B(DW5[0]), .Y(n3812) );
    znr8b U1007 ( .A(n3568), .B(DW6[29]), .C(DW6[27]), .D(DW6[30]), .E(DW6[23]
        ), .F(DW6[26]), .G(DW6[25]), .H(DW6[28]), .Y(n3567) );
    zor2b U1008 ( .A(QHSM[1]), .B(n3811), .Y(n3813) );
    zor2b U1009 ( .A(n3751), .B(n3749), .Y(n3750) );
    zivb U1010 ( .A(n3749), .Y(ACCEPT_DATA) );
    zoa211b U1011 ( .A(n3549), .B(n3129), .C(n2894), .D(n3551), .Y(n3550) );
    zoa211b U1012 ( .A(n3617), .B(n2920), .C(n3620), .D(n3621), .Y(n3619) );
    znr8b U1013 ( .A(VIR_TOTALBYTES_14), .B(VIR_TOTALBYTES_13), .C(n3618), .D(
        VIR_TOTALBYTES_9), .E(VIR_TOTALBYTES_12), .F(VIR_TOTALBYTES_7), .G(
        VIR_TOTALBYTES_1), .H(VIR_TOTALBYTES_0), .Y(n3617) );
    zivb U1014 ( .A(RXNAK), .Y(n3621) );
    zor2b U1015 ( .A(n3632), .B(n3840), .Y(n3841) );
    zmux21lb U1016 ( .A(n3623), .B(n3625), .S(n3774), .Y(n3840) );
    zoa22b U1017 ( .A(n2896), .B(n3570), .C(PCIEND), .D(n3571), .Y(n3569) );
    zan3b U1018 ( .A(DW6[7]), .B(n3488), .C(n3489), .Y(n3487) );
    zivb U1019 ( .A(SPD), .Y(n3786) );
    zivb U1020 ( .A(n3548), .Y(n3751) );
    zor2b U1021 ( .A(CERR_1), .B(n3773), .Y(n3624) );
    zivb U1022 ( .A(n3773), .Y(n3923) );
    zor2b U1023 ( .A(RXSTALL), .B(BABBLE), .Y(n3787) );
    zao32b U1024 ( .A(n3606), .B(n3133), .C(n3768), .D(n3766), .E(n3752), .Y(
        n3843) );
    zan2b U1025 ( .A(n3766), .B(n3620), .Y(n3842) );
    zor2b U1026 ( .A(n3753), .B(n3750), .Y(n3752) );
    zor2b U1027 ( .A(n3116), .B(n3596), .Y(n3605) );
    zor2b U1028 ( .A(n3516), .B(n2868), .Y(n3556) );
    zaoi2x4b U1029 ( .A(n2874), .B(n3591), .C(FEMPTY), .D(n3847), .E(n3848), 
        .F(n3105), .G(n3849), .H(n3497), .Y(n3524) );
    zoa22b U1030 ( .A(n3496), .B(n3497), .C(FEMPTY), .D(n3498), .Y(n3495) );
    zivb U1031 ( .A(n3496), .Y(n3849) );
    zivb U1032 ( .A(n3498), .Y(n3847) );
    zor2b U1033 ( .A(MULT_1), .B(MULT_0), .Y(n3626) );
    zor2b U1034 ( .A(QCMDSTART), .B(n3124), .Y(n3091) );
    zor2b U1035 ( .A(QHSM[6]), .B(QHSM[8]), .Y(n3532) );
    zivb U1036 ( .A(n3532), .Y(n3855) );
    zcx7b U1037 ( .A(TDMAEND), .B(n3126), .C(n3592), .D(n3595), .E(n3113), .Y(
        n3594) );
    znr6b U1038 ( .A(n3593), .B(MAXLEN[1]), .C(MAXLEN[0]), .D(MAXLEN[2]), .E(
        MAXLEN[4]), .F(MAXLEN[3]), .Y(n3592) );
    znd8b U1039 ( .A(n3685), .B(n3684), .C(n3682), .D(n3687), .E(n3686), .F(
        n3688), .G(n3683), .H(n3681), .Y(n3554) );
    zivb U1040 ( .A(DW2[3]), .Y(n3685) );
    zivc U1041 ( .A(DW2[1]), .Y(n3687) );
    zivb U1042 ( .A(DW2[2]), .Y(n3686) );
    zivc U1043 ( .A(DW2[7]), .Y(n3681) );
    zivd U1044 ( .A(n2919), .Y(n3329) );
    zor2b U1045 ( .A(n3100), .B(TRAN_CMD[14]), .Y(n3920) );
    zmux21lb U1046 ( .A(CPAGE_2), .B(CPAGE1177_2), .S(n2869), .Y(n3629) );
    zmux21lb U1047 ( .A(CPAGE_1), .B(CPAGE1177_1), .S(n2869), .Y(n3628) );
    zmux21lb U1048 ( .A(CPAGE_0), .B(n3739), .S(n2869), .Y(n3630) );
    zivb U1049 ( .A(CUROFFSET_T_12), .Y(n3743) );
    zaoi2x4b U1050 ( .A(DW10[0]), .B(n3866), .C(DW8[0]), .D(n3867), .E(DW9[0]), 
        .F(n3869), .G(DW5[0]), .H(n3868), .Y(n3905) );
    zao22b U1051 ( .A(DW9[1]), .B(n3869), .C(DW5[1]), .D(n3868), .Y(n3904) );
    zao22b U1052 ( .A(DW8[1]), .B(n3867), .C(DW10[1]), .D(n3866), .Y(n3903) );
    zao22b U1053 ( .A(DW9[2]), .B(n3869), .C(DW5[2]), .D(n3868), .Y(n3892) );
    zao22b U1054 ( .A(DW8[2]), .B(n3867), .C(DW10[2]), .D(n3866), .Y(n3891) );
    zao22b U1055 ( .A(DW9[3]), .B(n3869), .C(DW5[3]), .D(n3868), .Y(n3880) );
    zao22b U1056 ( .A(DW8[3]), .B(n3867), .C(DW10[3]), .D(n3866), .Y(n3879) );
    zao22b U1057 ( .A(DW9[4]), .B(n3869), .C(DW5[4]), .D(n3868), .Y(n3876) );
    zao22b U1058 ( .A(DW8[4]), .B(n3867), .C(DW10[4]), .D(n3866), .Y(n3875) );
    zaoi2x4b U1059 ( .A(DW10[5]), .B(n3866), .C(DW8[5]), .D(n3867), .E(DW5[5]), 
        .F(n3868), .G(n3869), .H(DW9[5]), .Y(n3873) );
    zaoi2x4b U1060 ( .A(DW10[6]), .B(n3866), .C(DW8[6]), .D(n3867), .E(DW5[6]), 
        .F(n3868), .G(n3869), .H(DW9[6]), .Y(n3872) );
    zaoi2x4b U1061 ( .A(DW10[7]), .B(n3866), .C(DW8[7]), .D(n3867), .E(DW5[7]), 
        .F(n3868), .G(n3869), .H(DW9[7]), .Y(n3871) );
    zaoi2x4b U1062 ( .A(DW10[8]), .B(n3866), .C(DW8[8]), .D(n3867), .E(DW5[8]), 
        .F(n3868), .G(n3869), .H(DW9[8]), .Y(n3870) );
    zaoi2x4b U1063 ( .A(n3866), .B(DW10[9]), .C(n3867), .D(DW8[9]), .E(n3868), 
        .F(DW5[9]), .G(n3869), .H(DW9[9]), .Y(n3862) );
    zaoi2x4b U1064 ( .A(DW10[10]), .B(n3866), .C(DW8[10]), .D(n3867), .E(DW5
        [10]), .F(n3868), .G(n3869), .H(DW9[10]), .Y(n3902) );
    zaoi2x4b U1065 ( .A(DW10[11]), .B(n3866), .C(DW8[11]), .D(n3867), .E(DW5
        [11]), .F(n3868), .G(n3869), .H(DW9[11]), .Y(n3901) );
    zoai2x4b U1066 ( .A(n3950), .B(n3222), .C(n3404), .D(n3802), .E(n3406), 
        .F(n3804), .G(n3408), .H(n3801), .Y(n3900) );
    zoai2x4b U1067 ( .A(n3949), .B(n3218), .C(n3411), .D(n3952), .E(n3412), 
        .F(n3954), .G(n3413), .H(n3956), .Y(n3899) );
    zoai2x4b U1068 ( .A(n3950), .B(n3210), .C(n3419), .D(n3952), .E(n3420), 
        .F(n3804), .G(n3421), .H(n3801), .Y(n3897) );
    zoai2x4b U1069 ( .A(n3949), .B(n3206), .C(n3423), .D(n3951), .E(n3424), 
        .F(n3954), .G(n3425), .H(n3955), .Y(n3896) );
    zoai2x4b U1070 ( .A(n3803), .B(n3202), .C(n3427), .D(n3802), .E(n3428), 
        .F(n3953), .G(n3429), .H(n3956), .Y(n3895) );
    zoai2x4b U1071 ( .A(n3950), .B(n3198), .C(n3431), .D(n3952), .E(n3432), 
        .F(n3804), .G(n3433), .H(n3801), .Y(n3894) );
    zoai2x4b U1072 ( .A(n3949), .B(n3194), .C(n3435), .D(n3951), .E(n3436), 
        .F(n3954), .G(n3437), .H(n3956), .Y(n3893) );
    zoai2x4b U1073 ( .A(n3803), .B(n3190), .C(n3439), .D(n3802), .E(n3440), 
        .F(n3953), .G(n3441), .H(n3955), .Y(n3890) );
    zoai2x4b U1074 ( .A(n3950), .B(n3186), .C(n3443), .D(n3952), .E(n3444), 
        .F(n3804), .G(n3445), .H(n3801), .Y(n3889) );
    zoai2x4b U1075 ( .A(n3949), .B(n3182), .C(n3447), .D(n3951), .E(n3448), 
        .F(n3954), .G(n3449), .H(n3956), .Y(n3888) );
    zoai2x4b U1076 ( .A(n3803), .B(n3178), .C(n3451), .D(n3802), .E(n3452), 
        .F(n3953), .G(n3453), .H(n3955), .Y(n3887) );
    zoai2x4b U1077 ( .A(n3950), .B(n3174), .C(n3455), .D(n3952), .E(n3456), 
        .F(n3804), .G(n3457), .H(n3801), .Y(n3886) );
    zoai2x4b U1078 ( .A(n3949), .B(n3170), .C(n3459), .D(n3951), .E(n3460), 
        .F(n3954), .G(n3461), .H(n3956), .Y(n3885) );
    zoai2x4b U1079 ( .A(n3803), .B(n3166), .C(n3463), .D(n3802), .E(n3464), 
        .F(n3953), .G(n3465), .H(n3955), .Y(n3884) );
    zoai2x4b U1080 ( .A(n3950), .B(n3162), .C(n3467), .D(n3952), .E(n3468), 
        .F(n3804), .G(n3469), .H(n3801), .Y(n3883) );
    zoai2x4b U1081 ( .A(n3949), .B(n3158), .C(n3471), .D(n3951), .E(n3472), 
        .F(n3954), .G(n3473), .H(n3956), .Y(n3882) );
    zivc U1082 ( .A(n3956), .Y(n3866) );
    zoai2x4b U1083 ( .A(n3803), .B(n3154), .C(n3475), .D(n3802), .E(n3476), 
        .F(n3953), .G(n3477), .H(n3955), .Y(n3881) );
    zivc U1084 ( .A(n3803), .Y(n3868) );
    zivc U1085 ( .A(n3802), .Y(n3867) );
    zivc U1086 ( .A(n3953), .Y(n3869) );
    zoai2x4b U1087 ( .A(n3950), .B(n3150), .C(n3479), .D(n3952), .E(n3480), 
        .F(n3804), .G(n3481), .H(n3801), .Y(n3878) );
    zor2b U1088 ( .A(n3794), .B(n3796), .Y(n3800) );
    zivb U1089 ( .A(DWCNT[3]), .Y(n3796) );
    zivb U1090 ( .A(n3798), .Y(n3919) );
    zor2b U1091 ( .A(DWCNT[0]), .B(DWCNT[3]), .Y(n3798) );
    zivb U1092 ( .A(n3791), .Y(n3908) );
    zoai2x4b U1093 ( .A(n3949), .B(n3145), .C(n3483), .D(n3951), .E(n3484), 
        .F(n3954), .G(n3485), .H(n3955), .Y(n3877) );
    zor2b U1094 ( .A(DWCNT[3]), .B(n3794), .Y(n3795) );
    zivb U1095 ( .A(DWCNT[0]), .Y(n3789) );
    znd2b U1096 ( .A(DW1[7]), .B(TRAN_CMD[6]), .Y(n3644) );
    zoai2x4b U1097 ( .A(PCIEND), .B(n3782), .C(n3565), .D(n3643), .E(n3493), 
        .F(n3784), .G(n3561), .H(n3588), .Y(n3906) );
    zivb U1098 ( .A(n3581), .Y(n3562) );
    zor2b U1099 ( .A(QHSM[4]), .B(QHSM[1]), .Y(n3586) );
    zan2b U1100 ( .A(n3580), .B(n3581), .Y(n3579) );
    zivb U1101 ( .A(n3563), .Y(n3580) );
    zivb U1102 ( .A(n3564), .Y(n3587) );
    zmux21lb U1103 ( .A(n3836), .B(n3582), .S(QHSM[2]), .Y(n3835) );
    zivb U1104 ( .A(n3644), .Y(n3577) );
    zmux21lb U1105 ( .A(n2876), .B(n3622), .S(PCIEND), .Y(n3834) );
    zan3b U1106 ( .A(n3575), .B(n3590), .C(n3493), .Y(n3622) );
    zivb U1107 ( .A(n3782), .Y(n3575) );
    zmux21lb U1108 ( .A(n3611), .B(n3740), .S(n3327), .Y(CERR1251_1) );
    zan2b U1109 ( .A(n3612), .B(n3613), .Y(n3611) );
    zmux21lb U1110 ( .A(n3614), .B(n3741), .S(LDPARM), .Y(CERR1251_0) );
    zan2b U1111 ( .A(n3615), .B(n3613), .Y(n3614) );
    zmux31hb U1112 ( .A(n2870), .B(n3327), .D0(MULT_1), .D1(MULT572_1), .D2(
        n3837), .Y(MULT588_1) );
    zxo2b U1113 ( .A(n3029), .B(MULT_0), .Y(MULT572_1) );
    zan3b U1114 ( .A(DW2[31]), .B(n3100), .C(n3554), .Y(n3837) );
    zmux31hb U1115 ( .A(n2870), .B(LDPARM), .D0(MULT_0), .D1(MULT572_0), .D2(
        n3838), .Y(MULT588_0) );
    zivb U1116 ( .A(n3626), .Y(n3642) );
    zivb U1117 ( .A(VIR_TOTALBYTES_11), .Y(n3762) );
    zivb U1118 ( .A(MINUEND_10), .Y(sub_457_B_not_10) );
    zivb U1119 ( .A(VIR_TOTALBYTES_10), .Y(n3763) );
    zivb U1120 ( .A(MINUEND_9), .Y(sub_457_B_not_9) );
    zivb U1121 ( .A(MINUEND_8), .Y(sub_457_B_not_8) );
    zivb U1122 ( .A(VIR_TOTALBYTES_8), .Y(n3756) );
    zivb U1123 ( .A(MINUEND_7), .Y(sub_457_B_not_7) );
    zivb U1124 ( .A(MINUEND_6), .Y(sub_457_B_not_6) );
    zivb U1125 ( .A(VIR_TOTALBYTES_6), .Y(n3757) );
    zivb U1126 ( .A(MINUEND_5), .Y(sub_457_B_not_5) );
    zivb U1127 ( .A(VIR_TOTALBYTES_5), .Y(n3758) );
    zivb U1128 ( .A(MINUEND_4), .Y(sub_457_B_not_4) );
    zivb U1129 ( .A(VIR_TOTALBYTES_4), .Y(n3759) );
    zivb U1130 ( .A(MINUEND_3), .Y(sub_457_B_not_3) );
    zivb U1131 ( .A(VIR_TOTALBYTES_3), .Y(n3760) );
    zivb U1132 ( .A(VIR_TOTALBYTES_2), .Y(n3761) );
    zivd U1133 ( .A(n3755), .Y(n3326) );
    zor2b U1134 ( .A(n3327), .B(n3620), .Y(n3755) );
    zivb U1135 ( .A(n3752), .Y(n3620) );
    zivd U1136 ( .A(n3754), .Y(n3328) );
    zor2b U1137 ( .A(n2920), .B(n3752), .Y(n3754) );
    zxo3b add_508_U1_6 ( .A(ACTLEN[6]), .B(UP_DW9[11]), .C(add_508_carry_6), 
        .Y(SBYTES966_6) );
    zivb U1138 ( .A(n3770), .Y(n3769) );
    zivf U1139 ( .A(n3765), .Y(n3322) );
    zivb U1140 ( .A(n3772), .Y(n3323) );
    zxo2b U1141 ( .A(r489_carry_2), .B(CPAGE_2), .Y(CPAGE1177_2) );
    zivb U1142 ( .A(n3818), .Y(n3817) );
    zhadrb r489_U1_1_1 ( .A(CPAGE_1), .B(CPAGE_0), .CO(r489_carry_2), .S(
        CPAGE1177_1) );
    zivf U1143 ( .A(FRNUM[2]), .Y(n3657) );
    zivf U1144 ( .A(FRNUM[1]), .Y(n3656) );
    zivf U1145 ( .A(FRNUM[0]), .Y(n3655) );
    zivb U1146 ( .A(n3605), .Y(n3768) );
    zivf U1147 ( .A(n3816), .Y(n3345) );
    zao2x4b U1148 ( .A(n2872), .B(UP_DW9[4]), .C(DW9[4]), .D(QH_PARSE_GO), .E(
        n3251), .F(FRNUM[7]), .G(FRAMETAG1498_4), .H(n2883), .Y(FRAMETAG1470_4
        ) );
    zxo2b U1149 ( .A(r469_carry_4), .B(FRNUM[7]), .Y(FRAMETAG1498_4) );
    zao2x4b U1150 ( .A(n2872), .B(UP_DW9[3]), .C(DW9[3]), .D(QH_PARSE_GO), .E(
        n3251), .F(FRNUM[6]), .G(FRAMETAG1498_3), .H(n2883), .Y(FRAMETAG1470_3
        ) );
    zhadrb r469_U1_1_3 ( .A(FRNUM[6]), .B(r469_carry_3), .CO(r469_carry_4), 
        .S(FRAMETAG1498_3) );
    zao2x4b U1151 ( .A(n2872), .B(UP_DW9[2]), .C(DW9[2]), .D(QH_PARSE_GO), .E(
        n3251), .F(FRNUM[5]), .G(FRAMETAG1498_2), .H(n2883), .Y(FRAMETAG1470_2
        ) );
    zhadrb r469_U1_1_2 ( .A(FRNUM[5]), .B(r469_carry_2), .CO(r469_carry_3), 
        .S(FRAMETAG1498_2) );
    zao2x4b U1152 ( .A(n2872), .B(UP_DW9[1]), .C(DW9[1]), .D(QH_PARSE_GO), .E(
        n3251), .F(FRNUM[4]), .G(FRAMETAG1498_1), .H(n2883), .Y(FRAMETAG1470_1
        ) );
    zivf U1153 ( .A(n3603), .Y(n3354) );
    zhadrb r469_U1_1_1 ( .A(FRNUM[4]), .B(FRNUM[3]), .CO(r469_carry_2), .S(
        FRAMETAG1498_1) );
    zao2x4b U1154 ( .A(n2872), .B(UP_DW9[0]), .C(DW9[0]), .D(QH_PARSE_GO), .E(
        n3251), .F(FRNUM[3]), .G(FRAMETAG1498_0), .H(n2883), .Y(FRAMETAG1470_0
        ) );
    zivb U1155 ( .A(n3767), .Y(n3810) );
    zivf U1156 ( .A(n3808), .Y(n3251) );
    zivb U1157 ( .A(n3604), .Y(n3809) );
    zivb U1158 ( .A(FRNUM[3]), .Y(FRAMETAG1498_0) );
    zoai2x4b U1159 ( .A(n3139), .B(n3927), .C(n3141), .D(n3142), .E(n3143), 
        .F(n3929), .G(n3145), .H(n3931), .Y(CURQTDPTR1736_31) );
    zivb U1160 ( .A(DW3[31]), .Y(n3139) );
    zivb U1161 ( .A(DW4[31]), .Y(n3143) );
    zivb U1162 ( .A(DW5[31]), .Y(n3145) );
    zoai2x4b U1163 ( .A(n3147), .B(n3926), .C(n3928), .D(n3148), .E(n3149), 
        .F(n3930), .G(n3150), .H(n3932), .Y(CURQTDPTR1736_30) );
    zivb U1164 ( .A(DW3[30]), .Y(n3147) );
    zivb U1165 ( .A(DW4[30]), .Y(n3149) );
    zivb U1166 ( .A(DW5[30]), .Y(n3150) );
    zivb U1167 ( .A(DW3[29]), .Y(n3151) );
    zivb U1168 ( .A(DW4[29]), .Y(n3153) );
    zivb U1169 ( .A(DW5[29]), .Y(n3154) );
    zoai2x4b U1170 ( .A(n3155), .B(n3927), .C(n3928), .D(n3156), .E(n3157), 
        .F(n3929), .G(n3158), .H(n3931), .Y(CURQTDPTR1736_28) );
    zivb U1171 ( .A(DW3[28]), .Y(n3155) );
    zivb U1172 ( .A(DW4[28]), .Y(n3157) );
    zivb U1173 ( .A(DW5[28]), .Y(n3158) );
    zoai2x4b U1174 ( .A(n3159), .B(n3926), .C(n3141), .D(n3160), .E(n3161), 
        .F(n3930), .G(n3162), .H(n3932), .Y(CURQTDPTR1736_27) );
    zivb U1175 ( .A(DW3[27]), .Y(n3159) );
    zivb U1176 ( .A(DW4[27]), .Y(n3161) );
    zivb U1177 ( .A(DW5[27]), .Y(n3162) );
    zivb U1178 ( .A(DW3[26]), .Y(n3163) );
    zivb U1179 ( .A(DW4[26]), .Y(n3165) );
    zivb U1180 ( .A(DW5[26]), .Y(n3166) );
    zivb U1181 ( .A(DW3[25]), .Y(n3167) );
    zivb U1182 ( .A(DW4[25]), .Y(n3169) );
    zivb U1183 ( .A(DW5[25]), .Y(n3170) );
    zoai2x4b U1184 ( .A(n3171), .B(n3926), .C(n3141), .D(n3172), .E(n3173), 
        .F(n3930), .G(n3174), .H(n3932), .Y(CURQTDPTR1736_24) );
    zivb U1185 ( .A(DW3[24]), .Y(n3171) );
    zivb U1186 ( .A(DW4[24]), .Y(n3173) );
    zivb U1187 ( .A(DW5[24]), .Y(n3174) );
    zivb U1188 ( .A(DW3[23]), .Y(n3175) );
    zivb U1189 ( .A(DW4[23]), .Y(n3177) );
    zivb U1190 ( .A(DW5[23]), .Y(n3178) );
    zoai2x4b U1191 ( .A(n3179), .B(n3926), .C(n3141), .D(n3180), .E(n3181), 
        .F(n3929), .G(n3182), .H(n3931), .Y(CURQTDPTR1736_22) );
    zivb U1192 ( .A(DW3[22]), .Y(n3179) );
    zivb U1193 ( .A(DW4[22]), .Y(n3181) );
    zivb U1194 ( .A(DW5[22]), .Y(n3182) );
    zivb U1195 ( .A(DW3[21]), .Y(n3183) );
    zivb U1196 ( .A(DW4[21]), .Y(n3185) );
    zivb U1197 ( .A(DW5[21]), .Y(n3186) );
    zoai2x4b U1198 ( .A(n3187), .B(n3140), .C(n3928), .D(n3188), .E(n3189), 
        .F(n3144), .G(n3190), .H(n3146), .Y(CURQTDPTR1736_20) );
    zivb U1199 ( .A(DW3[20]), .Y(n3187) );
    zivb U1200 ( .A(DW4[20]), .Y(n3189) );
    zivb U1201 ( .A(DW5[20]), .Y(n3190) );
    zoai2x4b U1202 ( .A(n3191), .B(n3926), .C(n3141), .D(n3192), .E(n3193), 
        .F(n3929), .G(n3194), .H(n3931), .Y(CURQTDPTR1736_19) );
    zivb U1203 ( .A(DW3[19]), .Y(n3191) );
    zivb U1204 ( .A(DW4[19]), .Y(n3193) );
    zivb U1205 ( .A(DW5[19]), .Y(n3194) );
    zivb U1206 ( .A(DW3[18]), .Y(n3195) );
    zivb U1207 ( .A(DW4[18]), .Y(n3197) );
    zivb U1208 ( .A(DW5[18]), .Y(n3198) );
    zivb U1209 ( .A(DW3[17]), .Y(n3199) );
    zivb U1210 ( .A(DW4[17]), .Y(n3201) );
    zivb U1211 ( .A(DW5[17]), .Y(n3202) );
    zoai2x4b U1212 ( .A(n3203), .B(n3926), .C(n3928), .D(n3204), .E(n3205), 
        .F(n3929), .G(n3206), .H(n3931), .Y(CURQTDPTR1736_16) );
    zivb U1213 ( .A(DW3[16]), .Y(n3203) );
    zivb U1214 ( .A(DW4[16]), .Y(n3205) );
    zivb U1215 ( .A(DW5[16]), .Y(n3206) );
    zoai2x4b U1216 ( .A(n3207), .B(n3927), .C(n3141), .D(n3208), .E(n3209), 
        .F(n3930), .G(n3210), .H(n3932), .Y(CURQTDPTR1736_15) );
    zivb U1217 ( .A(DW3[15]), .Y(n3207) );
    zivb U1218 ( .A(DW4[15]), .Y(n3209) );
    zivb U1219 ( .A(DW5[15]), .Y(n3210) );
    zivb U1220 ( .A(DW3[14]), .Y(n3211) );
    zivb U1221 ( .A(DW4[14]), .Y(n3213) );
    zivb U1222 ( .A(DW5[14]), .Y(n3214) );
    zoai2x4b U1223 ( .A(n3215), .B(n3926), .C(n3141), .D(n3216), .E(n3217), 
        .F(n3929), .G(n3218), .H(n3931), .Y(CURQTDPTR1736_13) );
    zivb U1224 ( .A(DW3[13]), .Y(n3215) );
    zivb U1225 ( .A(DW4[13]), .Y(n3217) );
    zivb U1226 ( .A(DW5[13]), .Y(n3218) );
    zivb U1227 ( .A(DW3[12]), .Y(n3219) );
    zivb U1228 ( .A(DW4[12]), .Y(n3221) );
    zivb U1229 ( .A(DW5[12]), .Y(n3222) );
    zivb U1230 ( .A(DW3[11]), .Y(n3223) );
    zivb U1231 ( .A(DW5[11]), .Y(n3226) );
    zoai2x4b U1232 ( .A(n3227), .B(n3926), .C(n3928), .D(n3228), .E(n3229), 
        .F(n3929), .G(n3230), .H(n3932), .Y(CURQTDPTR1736_10) );
    zivb U1233 ( .A(DW3[10]), .Y(n3227) );
    zivb U1234 ( .A(DW5[10]), .Y(n3230) );
    zivb U1235 ( .A(DW3[9]), .Y(n3231) );
    zivb U1236 ( .A(DW5[9]), .Y(n3234) );
    zoai2x4b U1237 ( .A(n3235), .B(n3140), .C(n3928), .D(n3236), .E(n3237), 
        .F(n3144), .G(n3238), .H(n3146), .Y(CURQTDPTR1736_8) );
    zivb U1238 ( .A(DW3[8]), .Y(n3235) );
    zivb U1239 ( .A(DW5[8]), .Y(n3238) );
    zivb U1240 ( .A(DW3[7]), .Y(n3239) );
    zivb U1241 ( .A(DW5[7]), .Y(n3242) );
    zoai2x4b U1242 ( .A(n3243), .B(n3926), .C(n3928), .D(n3244), .E(n3245), 
        .F(n3930), .G(n3246), .H(n3931), .Y(CURQTDPTR1736_6) );
    zivb U1243 ( .A(DW3[6]), .Y(n3243) );
    zivb U1244 ( .A(DW5[6]), .Y(n3246) );
    zoai2x4b U1245 ( .A(n3247), .B(n3140), .C(n3141), .D(n3248), .E(n3249), 
        .F(n3144), .G(n3250), .H(n3146), .Y(CURQTDPTR1736_5) );
    zivb U1246 ( .A(DW3[5]), .Y(n3247) );
    zivd U1247 ( .A(n3925), .Y(n3141) );
    zor2b U1248 ( .A(n3127), .B(n3133), .Y(n3925) );
    zivb U1249 ( .A(n3812), .Y(n3814) );
    zivb U1250 ( .A(DW5[5]), .Y(n3250) );
    zivd U1251 ( .A(n3925), .Y(n3928) );
    zivc U1252 ( .A(n3597), .Y(n3330) );
    zivb U1253 ( .A(n3750), .Y(n3922) );
    zivc U1254 ( .A(n3806), .Y(n3332) );
    zor2b U1255 ( .A(n3750), .B(n3360), .Y(n3806) );
    zivd U1256 ( .A(n3805), .Y(n3609) );
    zivd U1257 ( .A(n3748), .Y(n3608) );
    zan2b U1258 ( .A(n3105), .B(n3127), .Y(HCI_PRESOF_T1608) );
    zoai21b U1259 ( .A(n3118), .B(n3120), .C(n3121), .Y(PARSEQHEND_PRE) );
    zor2b U1260 ( .A(HCI_PRESOF), .B(HCI_PRESOF_T), .Y(n3105) );
    zor2b U1261 ( .A(QHSM[5]), .B(QHSM[7]), .Y(n3106) );
    zdffqrb QHSM_reg_9 ( .CK(PCICLK), .D(QHSMNXT_9), .R(TRST_), .Q(QHSM[9]) );
    zan2b U1262 ( .A(n3591), .B(QHSM[6]), .Y(n3107) );
    zivb U1263 ( .A(n3091), .Y(n3591) );
    zivb U1264 ( .A(n3105), .Y(n3566) );
    zivb U1265 ( .A(n3106), .Y(n3856) );
    zmux31lb U1266 ( .A(n3103), .B(n3327), .D0(n3104), .D1(n3831), .D2(n3648), 
        .Y(SPLITXSTATE1341) );
    zmux21lb U1267 ( .A(NXTISSTSWB), .B(n3830), .S(TRAN_CMD[14]), .Y(n3831) );
    zmux21lb U1268 ( .A(n3844), .B(n3578), .S(n3327), .Y(ACTIVE_NXT) );
    zoai21b U1269 ( .A(n3359), .B(n3360), .C(n3361), .Y(PING_ERR1014) );
    zivb U1270 ( .A(RXPIDERR), .Y(n3359) );
    zmux21lb U1271 ( .A(DW6[0]), .B(PING_ERR), .S(n3766), .Y(n3361) );
    zan3b U1272 ( .A(n3127), .B(n3133), .C(n3134), .Y(IMMEDRETRY1571) );
    zmux21lb U1273 ( .A(n3841), .B(n3491), .S(n3753), .Y(n3134) );
    zivb U1274 ( .A(n3811), .Y(QHSMNXT_1) );
    zor2b U1275 ( .A(n3531), .B(QRXERR), .Y(n3129) );
    zivb U1276 ( .A(n3129), .Y(n3774) );
    zmux21lb U1277 ( .A(n3534), .B(n3701), .S(n3327), .Y(XACTERR1308) );
    zan2b U1278 ( .A(n3535), .B(n3536), .Y(n3534) );
    zivb U1279 ( .A(PCIEND), .Y(n3116) );
    zoa211b U1280 ( .A(CACHE_INVALID), .B(n3133), .C(n3616), .D(n3596), .Y(
        n3119) );
    zor2b U1281 ( .A(n3097), .B(n3098), .Y(QHSMNXT_3) );
    zivb U1282 ( .A(n3643), .Y(n3490) );
    zoa211b U1283 ( .A(n3487), .B(n3492), .C(n3493), .D(n3090), .Y(n3098) );
    zivb U1284 ( .A(n3784), .Y(n3492) );
    zan2b U1285 ( .A(n3317), .B(n3133), .Y(CACHE_MODIFY502) );
    zmux21lb U1286 ( .A(n3599), .B(n3725), .S(LDPARM), .Y(MISUF1318) );
    zivb U1287 ( .A(n3556), .Y(n3522) );
    zoai21b U1288 ( .A(LTINT_PCLK), .B(n3135), .C(n3136), .Y(QHIOCINT_T2339)
         );
    zivb U1289 ( .A(EHCI_MAC_EOT), .Y(n3124) );
    zmux21lb U1290 ( .A(n3104), .B(n3764), .S(n3753), .Y(SPLITXSTATE_OLD1378)
         );
    zmux21lb U1291 ( .A(n3839), .B(n3641), .S(n3753), .Y(LENGTMAX867) );
    zivc U1292 ( .A(NXTISSTSWB), .Y(n3753) );
    zao21b U1293 ( .A(QHSMNXT_10), .B(n3093), .C(n3094), .Y(NXTISSTSWB) );
    zoa211b U1294 ( .A(QHERRINT), .B(n3131), .C(ERRINT_EN), .D(n3132), .Y(
        QHERRINT2450) );
    znd2b U1295 ( .A(ERRINT), .B(LTINT_PCLK), .Y(n3132) );
    zoa211b U1296 ( .A(QHIOCINT), .B(n3137), .C(USBINT_EN), .D(n3138), .Y(
        QHIOCINT2376) );
    zor2b U1297 ( .A(n3589), .B(n2881), .Y(n3137) );
    znd2b U1298 ( .A(USBINT), .B(LTINT_PCLK), .Y(n3138) );
    zivb U1299 ( .A(n3137), .Y(n3136) );
    zoai21b U1300 ( .A(LTINT_PCLK), .B(n3320), .C(n3321), .Y(QHERRINT_T2413)
         );
    zivb U1301 ( .A(n3131), .Y(n3321) );
    zivb U1302 ( .A(n3624), .Y(n3788) );
    zivd U1303 ( .A(n3121), .Y(LDPARM) );
    zor2b U1304 ( .A(QHSM[11]), .B(n3700), .Y(n3121) );
    zivb U1305 ( .A(QHSMNXT_3), .Y(n3700) );
    zivd U1306 ( .A(n3121), .Y(n3327) );
    zoai21b U1307 ( .A(n3355), .B(n3356), .C(n3357), .Y(DT1086) );
    zivb U1308 ( .A(DW1[14]), .Y(n3606) );
    zivd U1309 ( .A(QH_PARSE_GO), .Y(n3133) );
    zmux21lb U1310 ( .A(n3842), .B(n3843), .S(DT), .Y(n3357) );
    zan3b U1311 ( .A(DW6[7]), .B(n3090), .C(n3318), .Y(QHSMNXT_2) );
    zao32b U1312 ( .A(n3489), .B(n3488), .C(INACT_COND), .D(n3909), .E(PCIEND), 
        .Y(n3318) );
    zivb U1313 ( .A(n3650), .Y(n3489) );
    zivb U1314 ( .A(n3571), .Y(n3909) );
    zan2b U1315 ( .A(QHERRINT_T), .B(LTINT_PCLK), .Y(QHERRINT_S) );
    zan2b U1316 ( .A(LTINT_PCLK), .B(QHIOCINT_T), .Y(QHIOCINT_S) );
    znd8b U1317 ( .A(n3108), .B(n3109), .C(n3110), .D(n3111), .E(n3112), .F(
        n3113), .G(n3114), .H(n3115), .Y(QTDEXE) );
    zivb U1318 ( .A(QHSMNXT_7), .Y(n3108) );
    zao32b U1319 ( .A(n2875), .B(n3095), .C(n2882), .D(n2884), .E(TRAN_CMD
        [104]), .Y(QHSMNXT_7) );
    zivb U1320 ( .A(QCMDSTART), .Y(n3095) );
    zivb U1321 ( .A(QHSMNXT_5), .Y(n3110) );
    zao32b U1322 ( .A(n2873), .B(n3095), .C(n2882), .D(n2884), .E(n3096), .Y(
        QHSMNXT_5) );
    zivb U1323 ( .A(QHSMNXT_8), .Y(n3112) );
    zao33b U1324 ( .A(n3092), .B(n3090), .C(n3091), .D(QCMDSTART), .E(n2875), 
        .F(n2882), .Y(QHSMNXT_8) );
    zivb U1325 ( .A(n3776), .Y(n3092) );
    zivb U1326 ( .A(PHASENXT_outcyc), .Y(n3113) );
    zao33b U1327 ( .A(n2874), .B(n3090), .C(n3091), .D(n2873), .E(QCMDSTART), 
        .F(n2882), .Y(PHASENXT_outcyc) );
    zivb U1328 ( .A(n3109), .Y(QHSMNXT_9) );
    zivb U1329 ( .A(n3111), .Y(QHSMNXT_4) );
    zivb U1330 ( .A(n3114), .Y(QHSMNXT_10) );
    zivb U1331 ( .A(n3115), .Y(PHASENXT_resultwb) );
    zan2b U1332 ( .A(n3101), .B(n3102), .Y(QCMDSTART_REQ) );
    zivb U1333 ( .A(n3130), .Y(QBUI_GO) );
    zor2b U1334 ( .A(QHSM[4]), .B(n3111), .Y(n3130) );
    zan2b U1335 ( .A(n3103), .B(n3104), .Y(TRAN_CMD[0]) );
    zivb U1336 ( .A(n3631), .Y(n3103) );
    zor2b U1337 ( .A(n3632), .B(n3100), .Y(n3631) );
    zivb U1338 ( .A(n3554), .Y(n3632) );
    zor2b U1339 ( .A(TRAN_CMD[7]), .B(n3099), .Y(TRAN_CMD[4]) );
    zivb U1340 ( .A(TRAN_CMD[4]), .Y(TRAN_CMD[3]) );
    zan2b U1341 ( .A(n3125), .B(n2921), .Y(TRAN_CMD[8]) );
    zivb U1342 ( .A(DW6[9]), .Y(n3125) );
    zan2b U1343 ( .A(n3319), .B(MAXLEN[0]), .Y(TRAN_CMD[40]) );
    zan2b U1344 ( .A(n3319), .B(MAXLEN[1]), .Y(TRAN_CMD[41]) );
    zan2b U1345 ( .A(n3319), .B(MAXLEN[2]), .Y(TRAN_CMD[42]) );
    zan2b U1346 ( .A(n3319), .B(MAXLEN[3]), .Y(TRAN_CMD[43]) );
    zan2b U1347 ( .A(n3319), .B(MAXLEN[4]), .Y(TRAN_CMD[44]) );
    zan2b U1348 ( .A(n3319), .B(MAXLEN[5]), .Y(TRAN_CMD[45]) );
    zan2b U1349 ( .A(n3319), .B(MAXLEN[6]), .Y(TRAN_CMD[46]) );
    zan2b U1350 ( .A(n3319), .B(MAXLEN[7]), .Y(TRAN_CMD[47]) );
    zan2b U1351 ( .A(n3319), .B(MAXLEN[8]), .Y(TRAN_CMD[48]) );
    zan2b U1352 ( .A(n3319), .B(MAXLEN[9]), .Y(TRAN_CMD[49]) );
    zan2b U1353 ( .A(n3319), .B(MAXLEN[10]), .Y(TRAN_CMD[50]) );
    zivb U1354 ( .A(n3920), .Y(n3530) );
    zoai2x4b U1355 ( .A(n3936), .B(n3404), .C(n3405), .D(n3406), .E(n3940), 
        .F(n3408), .G(n3409), .H(n3410), .Y(TRAN_CMD[52]) );
    zivb U1356 ( .A(DW8[12]), .Y(n3404) );
    zivb U1357 ( .A(DW9[12]), .Y(n3406) );
    zivb U1358 ( .A(DW10[12]), .Y(n3408) );
    zivb U1359 ( .A(DW11[12]), .Y(n3410) );
    zoai2x4b U1360 ( .A(n3403), .B(n3411), .C(n3937), .D(n3412), .E(n3407), 
        .F(n3413), .G(n3409), .H(n3414), .Y(TRAN_CMD[53]) );
    zivb U1361 ( .A(DW8[13]), .Y(n3411) );
    zivb U1362 ( .A(DW9[13]), .Y(n3412) );
    zivb U1363 ( .A(DW10[13]), .Y(n3413) );
    zivb U1364 ( .A(DW11[13]), .Y(n3414) );
    zoai2x4b U1365 ( .A(n3935), .B(n3415), .C(n3938), .D(n3416), .E(n3939), 
        .F(n3417), .G(n3409), .H(n3418), .Y(TRAN_CMD[54]) );
    zivb U1366 ( .A(DW8[14]), .Y(n3415) );
    zivb U1367 ( .A(DW9[14]), .Y(n3416) );
    zivb U1368 ( .A(DW10[14]), .Y(n3417) );
    zivb U1369 ( .A(DW11[14]), .Y(n3418) );
    zoai2x4b U1370 ( .A(n3936), .B(n3419), .C(n3405), .D(n3420), .E(n3940), 
        .F(n3421), .G(n3409), .H(n3422), .Y(TRAN_CMD[55]) );
    zivb U1371 ( .A(DW8[15]), .Y(n3419) );
    zivb U1372 ( .A(DW9[15]), .Y(n3420) );
    zivb U1373 ( .A(DW10[15]), .Y(n3421) );
    zivb U1374 ( .A(DW11[15]), .Y(n3422) );
    zoai2x4b U1375 ( .A(n3403), .B(n3423), .C(n3938), .D(n3424), .E(n3407), 
        .F(n3425), .G(n3409), .H(n3426), .Y(TRAN_CMD[56]) );
    zivb U1376 ( .A(DW8[16]), .Y(n3423) );
    zivb U1377 ( .A(DW9[16]), .Y(n3424) );
    zivb U1378 ( .A(DW10[16]), .Y(n3425) );
    zivb U1379 ( .A(DW11[16]), .Y(n3426) );
    zoai2x4b U1380 ( .A(n3935), .B(n3427), .C(n3937), .D(n3428), .E(n3939), 
        .F(n3429), .G(n3409), .H(n3430), .Y(TRAN_CMD[57]) );
    zivb U1381 ( .A(DW8[17]), .Y(n3427) );
    zivb U1382 ( .A(DW9[17]), .Y(n3428) );
    zivb U1383 ( .A(DW10[17]), .Y(n3429) );
    zivb U1384 ( .A(DW11[17]), .Y(n3430) );
    zoai2x4b U1385 ( .A(n3936), .B(n3431), .C(n3405), .D(n3432), .E(n3940), 
        .F(n3433), .G(n3409), .H(n3434), .Y(TRAN_CMD[58]) );
    zivb U1386 ( .A(DW8[18]), .Y(n3431) );
    zivb U1387 ( .A(DW9[18]), .Y(n3432) );
    zivb U1388 ( .A(DW10[18]), .Y(n3433) );
    zivb U1389 ( .A(DW11[18]), .Y(n3434) );
    zoai2x4b U1390 ( .A(n3403), .B(n3435), .C(n3937), .D(n3436), .E(n3407), 
        .F(n3437), .G(n3409), .H(n3438), .Y(TRAN_CMD[59]) );
    zivb U1391 ( .A(DW8[19]), .Y(n3435) );
    zivb U1392 ( .A(DW9[19]), .Y(n3436) );
    zivb U1393 ( .A(DW10[19]), .Y(n3437) );
    zivb U1394 ( .A(DW11[19]), .Y(n3438) );
    zoai2x4b U1395 ( .A(n3935), .B(n3439), .C(n3938), .D(n3440), .E(n3939), 
        .F(n3441), .G(n3409), .H(n3442), .Y(TRAN_CMD[60]) );
    zivb U1396 ( .A(DW8[20]), .Y(n3439) );
    zivb U1397 ( .A(DW9[20]), .Y(n3440) );
    zivb U1398 ( .A(DW10[20]), .Y(n3441) );
    zivb U1399 ( .A(DW11[20]), .Y(n3442) );
    zoai2x4b U1400 ( .A(n3936), .B(n3443), .C(n3405), .D(n3444), .E(n3940), 
        .F(n3445), .G(n3409), .H(n3446), .Y(TRAN_CMD[61]) );
    zivb U1401 ( .A(DW8[21]), .Y(n3443) );
    zivb U1402 ( .A(DW9[21]), .Y(n3444) );
    zivb U1403 ( .A(DW10[21]), .Y(n3445) );
    zivb U1404 ( .A(DW11[21]), .Y(n3446) );
    zoai2x4b U1405 ( .A(n3403), .B(n3447), .C(n3938), .D(n3448), .E(n3407), 
        .F(n3449), .G(n3409), .H(n3450), .Y(TRAN_CMD[62]) );
    zivb U1406 ( .A(DW8[22]), .Y(n3447) );
    zivb U1407 ( .A(DW9[22]), .Y(n3448) );
    zivb U1408 ( .A(DW10[22]), .Y(n3449) );
    zivb U1409 ( .A(DW11[22]), .Y(n3450) );
    zoai2x4b U1410 ( .A(n3935), .B(n3451), .C(n3405), .D(n3452), .E(n3939), 
        .F(n3453), .G(n3409), .H(n3454), .Y(TRAN_CMD[63]) );
    zivb U1411 ( .A(DW8[23]), .Y(n3451) );
    zivb U1412 ( .A(DW9[23]), .Y(n3452) );
    zivb U1413 ( .A(DW10[23]), .Y(n3453) );
    zivb U1414 ( .A(DW11[23]), .Y(n3454) );
    zoai2x4b U1415 ( .A(n3936), .B(n3455), .C(n3937), .D(n3456), .E(n3940), 
        .F(n3457), .G(n3409), .H(n3458), .Y(TRAN_CMD[64]) );
    zivb U1416 ( .A(DW8[24]), .Y(n3455) );
    zivb U1417 ( .A(DW9[24]), .Y(n3456) );
    zivb U1418 ( .A(DW10[24]), .Y(n3457) );
    zivb U1419 ( .A(DW11[24]), .Y(n3458) );
    zoai2x4b U1420 ( .A(n3403), .B(n3459), .C(n3937), .D(n3460), .E(n3407), 
        .F(n3461), .G(n3409), .H(n3462), .Y(TRAN_CMD[65]) );
    zivb U1421 ( .A(DW8[25]), .Y(n3459) );
    zivb U1422 ( .A(DW9[25]), .Y(n3460) );
    zivb U1423 ( .A(DW10[25]), .Y(n3461) );
    zivb U1424 ( .A(DW11[25]), .Y(n3462) );
    zoai2x4b U1425 ( .A(n3935), .B(n3463), .C(n3938), .D(n3464), .E(n3939), 
        .F(n3465), .G(n3409), .H(n3466), .Y(TRAN_CMD[66]) );
    zivb U1426 ( .A(DW8[26]), .Y(n3463) );
    zivb U1427 ( .A(DW9[26]), .Y(n3464) );
    zivb U1428 ( .A(DW10[26]), .Y(n3465) );
    zivb U1429 ( .A(DW11[26]), .Y(n3466) );
    zoai2x4b U1430 ( .A(n3467), .B(n3935), .C(n3468), .D(n3937), .E(n3469), 
        .F(n3407), .G(n3409), .H(n3470), .Y(TRAN_CMD[67]) );
    zivb U1431 ( .A(DW8[27]), .Y(n3467) );
    zivb U1432 ( .A(DW9[27]), .Y(n3468) );
    zivb U1433 ( .A(DW10[27]), .Y(n3469) );
    zivb U1434 ( .A(DW11[27]), .Y(n3470) );
    zoai2x4b U1435 ( .A(n3936), .B(n3471), .C(n3405), .D(n3472), .E(n3940), 
        .F(n3473), .G(n3409), .H(n3474), .Y(TRAN_CMD[68]) );
    zivb U1436 ( .A(DW8[28]), .Y(n3471) );
    zivb U1437 ( .A(DW9[28]), .Y(n3472) );
    zivb U1438 ( .A(DW10[28]), .Y(n3473) );
    zivb U1439 ( .A(DW11[28]), .Y(n3474) );
    zoai2x4b U1440 ( .A(n3403), .B(n3475), .C(n3937), .D(n3476), .E(n3407), 
        .F(n3477), .G(n3409), .H(n3478), .Y(TRAN_CMD[69]) );
    zivb U1441 ( .A(DW8[29]), .Y(n3475) );
    zivb U1442 ( .A(DW9[29]), .Y(n3476) );
    zivb U1443 ( .A(DW10[29]), .Y(n3477) );
    zivb U1444 ( .A(DW11[29]), .Y(n3478) );
    zoai2x4b U1445 ( .A(n3935), .B(n3479), .C(n3938), .D(n3480), .E(n3939), 
        .F(n3481), .G(n3409), .H(n3482), .Y(TRAN_CMD[70]) );
    zivb U1446 ( .A(DW8[30]), .Y(n3479) );
    zivb U1447 ( .A(DW9[30]), .Y(n3480) );
    zivb U1448 ( .A(DW10[30]), .Y(n3481) );
    zivb U1449 ( .A(DW11[30]), .Y(n3482) );
    zoai2x4b U1450 ( .A(n3936), .B(n3483), .C(n3405), .D(n3484), .E(n3940), 
        .F(n3485), .G(n3409), .H(n3486), .Y(TRAN_CMD[71]) );
    zivb U1451 ( .A(DW8[31]), .Y(n3483) );
    zivb U1452 ( .A(DW9[31]), .Y(n3484) );
    zivb U1453 ( .A(DW10[31]), .Y(n3485) );
    zivf U1454 ( .A(n3921), .Y(n3409) );
    zao21b U1455 ( .A(n3746), .B(n3747), .C(n3745), .Y(n3921) );
    zivb U1456 ( .A(DW11[31]), .Y(n3486) );
    zan2b U1457 ( .A(DW8[12]), .B(n3543), .Y(n3401) );
    zan2b U1458 ( .A(DW8[13]), .B(n3543), .Y(n3399) );
    zan2b U1459 ( .A(DW8[14]), .B(n3543), .Y(n3397) );
    zan2b U1460 ( .A(DW8[15]), .B(n3543), .Y(n3395) );
    zan2b U1461 ( .A(DW8[16]), .B(n3543), .Y(n3393) );
    zan2b U1462 ( .A(DW8[17]), .B(n3543), .Y(n3391) );
    zan2b U1463 ( .A(DW8[18]), .B(n3543), .Y(n3389) );
    zan2b U1464 ( .A(DW8[19]), .B(n3543), .Y(n3387) );
    zan2b U1465 ( .A(DW8[20]), .B(n3543), .Y(n3385) );
    zan2b U1466 ( .A(DW8[21]), .B(n3543), .Y(n3383) );
    zan2b U1467 ( .A(DW8[22]), .B(n3543), .Y(n3381) );
    zan2b U1468 ( .A(DW8[23]), .B(n3543), .Y(n3379) );
    zan2b U1469 ( .A(DW8[24]), .B(n3543), .Y(n3377) );
    zan2b U1470 ( .A(DW8[25]), .B(n3543), .Y(n3375) );
    zan2b U1471 ( .A(DW8[26]), .B(n3543), .Y(n3373) );
    zan2b U1472 ( .A(n3543), .B(DW8[27]), .Y(n3371) );
    zan2b U1473 ( .A(DW8[28]), .B(n3543), .Y(n3369) );
    zan2b U1474 ( .A(DW8[29]), .B(n3543), .Y(n3367) );
    zan2b U1475 ( .A(DW8[30]), .B(n3543), .Y(n3365) );
    zivf U1476 ( .A(n3403), .Y(n3362) );
    zivb U1477 ( .A(n3630), .Y(n3746) );
    zivb U1478 ( .A(n3628), .Y(n3747) );
    zivd U1479 ( .A(n3629), .Y(n3745) );
    zan2b U1480 ( .A(DW8[31]), .B(n3543), .Y(n3363) );
    zivf U1481 ( .A(n3938), .Y(n3543) );
    zivd U1482 ( .A(n3629), .Y(n3948) );
    zivf U1483 ( .A(n3744), .Y(n3851) );
    zivf U1484 ( .A(n3939), .Y(n3852) );
    zivb U1485 ( .A(n3520), .Y(n3126) );
    zor2b U1486 ( .A(n3100), .B(n3104), .Y(n3520) );
    zivc U1487 ( .A(TRAN_CMD[6]), .Y(n3100) );
    zivb U1488 ( .A(TRAN_CMD[104]), .Y(n3096) );
    zoai21b U1489 ( .A(n3785), .B(n3792), .C(n3905), .Y(n3253) );
    zivb U1490 ( .A(DW4[0]), .Y(n3785) );
    zoai21b U1491 ( .A(n3792), .B(n3249), .C(n3873), .Y(n3263) );
    zivb U1492 ( .A(DW4[5]), .Y(n3249) );
    zoai21b U1493 ( .A(n3792), .B(n3245), .C(n3872), .Y(n3265) );
    zivb U1494 ( .A(DW4[6]), .Y(n3245) );
    zoai21b U1495 ( .A(n3792), .B(n3241), .C(n3871), .Y(n3267) );
    zivb U1496 ( .A(DW4[7]), .Y(n3241) );
    zoai21b U1497 ( .A(n3792), .B(n3237), .C(n3870), .Y(n3269) );
    zivb U1498 ( .A(DW4[8]), .Y(n3237) );
    zoai21b U1499 ( .A(n3792), .B(n3233), .C(n3862), .Y(n3271) );
    zivb U1500 ( .A(DW4[9]), .Y(n3233) );
    zoai21b U1501 ( .A(n3792), .B(n3229), .C(n3902), .Y(n3273) );
    zivb U1502 ( .A(DW4[10]), .Y(n3229) );
    zoai21b U1503 ( .A(n3792), .B(n3225), .C(n3901), .Y(n3275) );
    zivb U1504 ( .A(DW4[11]), .Y(n3225) );
    zao21b U1505 ( .A(DW4[12]), .B(n3874), .C(n3900), .Y(n3277) );
    zivc U1506 ( .A(n3792), .Y(n3874) );
    zao21b U1507 ( .A(DW4[13]), .B(n3947), .C(n3899), .Y(n3279) );
    zivc U1508 ( .A(n3792), .Y(n3947) );
    zao21b U1509 ( .A(DW4[14]), .B(n3874), .C(n3898), .Y(n3281) );
    zao21b U1510 ( .A(DW4[15]), .B(n3947), .C(n3897), .Y(n3283) );
    zao21b U1511 ( .A(DW4[16]), .B(n3874), .C(n3896), .Y(n3285) );
    zao21b U1512 ( .A(DW4[17]), .B(n3947), .C(n3895), .Y(n3287) );
    zao21b U1513 ( .A(DW4[18]), .B(n3874), .C(n3894), .Y(n3289) );
    zao21b U1514 ( .A(DW4[19]), .B(n3947), .C(n3893), .Y(n3291) );
    zao21b U1515 ( .A(DW4[20]), .B(n3874), .C(n3890), .Y(n3293) );
    zao21b U1516 ( .A(DW4[21]), .B(n3947), .C(n3889), .Y(n3295) );
    zao21b U1517 ( .A(DW4[22]), .B(n3874), .C(n3888), .Y(n3297) );
    zao21b U1518 ( .A(DW4[23]), .B(n3947), .C(n3887), .Y(n3299) );
    zao21b U1519 ( .A(DW4[24]), .B(n3874), .C(n3886), .Y(n3301) );
    zao21b U1520 ( .A(DW4[25]), .B(n3947), .C(n3885), .Y(n3303) );
    zao21b U1521 ( .A(DW4[26]), .B(n3874), .C(n3884), .Y(n3305) );
    zao21b U1522 ( .A(DW4[27]), .B(n3947), .C(n3883), .Y(n3307) );
    zao21b U1523 ( .A(DW4[28]), .B(n3874), .C(n3882), .Y(n3309) );
    zao21b U1524 ( .A(DW4[29]), .B(n3947), .C(n3881), .Y(n3311) );
    zao21b U1525 ( .A(DW4[30]), .B(n3874), .C(n3878), .Y(n3313) );
    zivd U1526 ( .A(n3800), .Y(n3863) );
    zivb U1527 ( .A(n3790), .Y(n3918) );
    zivb U1528 ( .A(n3795), .Y(n3907) );
    zao21b U1529 ( .A(DW4[31]), .B(n3947), .C(n3877), .Y(n3315) );
    zivd U1530 ( .A(n3800), .Y(n3942) );
    zivb U1531 ( .A(n3117), .Y(QHCIADR[4]) );
    zor2b U1532 ( .A(QHDWNUM[0]), .B(n3493), .Y(n3117) );
    zmux21hb U1533 ( .A(UP_DW3[5]), .B(CACHE_ADDR[0]), .S(n2931), .Y(QHCIADR
        [5]) );
    zmux21hb U1534 ( .A(UP_DW3[6]), .B(CACHE_ADDR[1]), .S(n2931), .Y(QHCIADR
        [6]) );
    zmux21hb U1535 ( .A(UP_DW3[7]), .B(CACHE_ADDR[2]), .S(n2931), .Y(QHCIADR
        [7]) );
    zmux21hb U1536 ( .A(UP_DW3[8]), .B(CACHE_ADDR[3]), .S(n2931), .Y(QHCIADR
        [8]) );
    zmux21hb U1537 ( .A(UP_DW3[9]), .B(CACHE_ADDR[4]), .S(QHSM[12]), .Y(
        QHCIADR[9]) );
    zmux21hb U1538 ( .A(UP_DW3[10]), .B(CACHE_ADDR[5]), .S(n2931), .Y(QHCIADR
        [10]) );
    zmux21hb U1539 ( .A(UP_DW3[11]), .B(CACHE_ADDR[6]), .S(n2931), .Y(QHCIADR
        [11]) );
    zmux21hb U1540 ( .A(UP_DW3[12]), .B(CACHE_ADDR[7]), .S(n2931), .Y(QHCIADR
        [12]) );
    zmux21hb U1541 ( .A(UP_DW3[13]), .B(CACHE_ADDR[8]), .S(n2931), .Y(QHCIADR
        [13]) );
    zmux21hb U1542 ( .A(UP_DW3[14]), .B(CACHE_ADDR[9]), .S(QHSM[12]), .Y(
        QHCIADR[14]) );
    zmux21hb U1543 ( .A(UP_DW3[15]), .B(CACHE_ADDR[10]), .S(n2931), .Y(QHCIADR
        [15]) );
    zmux21hb U1544 ( .A(UP_DW3[16]), .B(CACHE_ADDR[11]), .S(QHSM[12]), .Y(
        QHCIADR[16]) );
    zmux21hb U1545 ( .A(UP_DW3[17]), .B(CACHE_ADDR[12]), .S(QHSM[12]), .Y(
        QHCIADR[17]) );
    zmux21hb U1546 ( .A(UP_DW3[18]), .B(CACHE_ADDR[13]), .S(QHSM[12]), .Y(
        QHCIADR[18]) );
    zmux21hb U1547 ( .A(UP_DW3[19]), .B(CACHE_ADDR[14]), .S(QHSM[12]), .Y(
        QHCIADR[19]) );
    zmux21hb U1548 ( .A(UP_DW3[20]), .B(CACHE_ADDR[15]), .S(QHSM[12]), .Y(
        QHCIADR[20]) );
    zmux21hb U1549 ( .A(UP_DW3[21]), .B(CACHE_ADDR[16]), .S(QHSM[12]), .Y(
        QHCIADR[21]) );
    zmux21hb U1550 ( .A(UP_DW3[22]), .B(CACHE_ADDR[17]), .S(n2931), .Y(QHCIADR
        [22]) );
    zmux21hb U1551 ( .A(UP_DW3[23]), .B(CACHE_ADDR[18]), .S(QHSM[12]), .Y(
        QHCIADR[23]) );
    zmux21hb U1552 ( .A(UP_DW3[24]), .B(CACHE_ADDR[19]), .S(n2931), .Y(QHCIADR
        [24]) );
    zmux21hb U1553 ( .A(UP_DW3[25]), .B(CACHE_ADDR[20]), .S(QHSM[12]), .Y(
        QHCIADR[25]) );
    zmux21hb U1554 ( .A(UP_DW3[26]), .B(CACHE_ADDR[21]), .S(n2931), .Y(QHCIADR
        [26]) );
    zmux21hb U1555 ( .A(UP_DW3[27]), .B(CACHE_ADDR[22]), .S(QHSM[12]), .Y(
        QHCIADR[27]) );
    zmux21hb U1556 ( .A(UP_DW3[28]), .B(CACHE_ADDR[23]), .S(n2931), .Y(QHCIADR
        [28]) );
    zmux21hb U1557 ( .A(UP_DW3[29]), .B(CACHE_ADDR[24]), .S(QHSM[12]), .Y(
        QHCIADR[29]) );
    zmux21hb U1558 ( .A(UP_DW3[30]), .B(CACHE_ADDR[25]), .S(n2931), .Y(QHCIADR
        [30]) );
    zmux21hb U1559 ( .A(UP_DW3[31]), .B(CACHE_ADDR[26]), .S(QHSM[12]), .Y(
        QHCIADR[31]) );
    zor2b U1560 ( .A(QHDWNUM[0]), .B(INACT_COND), .Y(n3797) );
    zor2b U1561 ( .A(QHSM[1]), .B(QHCIMWR), .Y(QHCIREQ) );
    zor2b U1562 ( .A(QHSM[11]), .B(QHSM[2]), .Y(CACHEPHASE) );
    zor2b U1563 ( .A(UP_LDW7), .B(UP_CACHE1), .Y(UP_LDW6) );
    zmux21lb U1564 ( .A(n3829), .B(n3742), .S(n3324), .Y(UP_DW6[0]) );
    zivb U1565 ( .A(DW6[0]), .Y(n3742) );
    zmux21lb U1566 ( .A(n3104), .B(n3648), .S(n3941), .Y(UP_DW6[1]) );
    zivb U1567 ( .A(DW6[1]), .Y(n3648) );
    zmux21lb U1568 ( .A(n3601), .B(n3725), .S(n3941), .Y(UP_DW6[2]) );
    zivb U1569 ( .A(DW6[2]), .Y(n3725) );
    zmux21lb U1570 ( .A(n3535), .B(n3701), .S(n3324), .Y(UP_DW6[3]) );
    zivb U1571 ( .A(DW6[3]), .Y(n3701) );
    zao21b U1572 ( .A(BABBLE), .B(n3325), .C(DW6[4]), .Y(UP_DW6[4]) );
    zan2b U1573 ( .A(DW6[5]), .B(n3941), .Y(UP_DW6[5]) );
    zmux21lb U1574 ( .A(n3827), .B(n3488), .S(n3324), .Y(UP_DW6[6]) );
    zivb U1575 ( .A(DW6[6]), .Y(n3488) );
    zmux21lb U1576 ( .A(n3590), .B(n3826), .S(n3941), .Y(UP_DW6[7]) );
    zor2b U1577 ( .A(INACT_COND), .B(n3578), .Y(n3826) );
    zivb U1578 ( .A(DW6[7]), .Y(n3578) );
    zmux21lb U1579 ( .A(n3828), .B(n3741), .S(n3324), .Y(UP_DW6[10]) );
    zivb U1580 ( .A(DW6[10]), .Y(n3741) );
    zmux21lb U1581 ( .A(n3085), .B(n3740), .S(n3941), .Y(UP_DW6[11]) );
    zivb U1582 ( .A(DW6[11]), .Y(n3740) );
    zmux21lb U1583 ( .A(n3739), .B(n3738), .S(n3324), .Y(UP_DW6[12]) );
    zivb U1584 ( .A(DW6[12]), .Y(n3738) );
    zmux21lb U1585 ( .A(n3737), .B(n3736), .S(n3941), .Y(UP_DW6[13]) );
    zivb U1586 ( .A(DW6[13]), .Y(n3736) );
    zmux21lb U1587 ( .A(n3735), .B(n3734), .S(n3324), .Y(UP_DW6[14]) );
    zivb U1588 ( .A(DW6[14]), .Y(n3734) );
    zmux21lb U1589 ( .A(n3733), .B(n3732), .S(n3941), .Y(UP_DW6[16]) );
    zivb U1590 ( .A(DW6[16]), .Y(n3732) );
    zmux21lb U1591 ( .A(n3731), .B(n3730), .S(n3324), .Y(UP_DW6[17]) );
    zivb U1592 ( .A(DW6[17]), .Y(n3730) );
    zmux21lb U1593 ( .A(n3729), .B(n3728), .S(n3941), .Y(UP_DW6[18]) );
    zivb U1594 ( .A(DW6[18]), .Y(n3728) );
    zmux21lb U1595 ( .A(n3727), .B(n3726), .S(n3324), .Y(UP_DW6[19]) );
    zivb U1596 ( .A(DW6[19]), .Y(n3726) );
    zmux21lb U1597 ( .A(n3724), .B(n3723), .S(n3324), .Y(UP_DW6[20]) );
    zivb U1598 ( .A(DW6[20]), .Y(n3723) );
    zmux21lb U1599 ( .A(n3722), .B(n3721), .S(n3941), .Y(UP_DW6[21]) );
    zivb U1600 ( .A(DW6[21]), .Y(n3721) );
    zmux21lb U1601 ( .A(n3720), .B(n3719), .S(n3324), .Y(UP_DW6[22]) );
    zivb U1602 ( .A(DW6[22]), .Y(n3719) );
    zmux21lb U1603 ( .A(n3718), .B(n3717), .S(n3941), .Y(UP_DW6[23]) );
    zivb U1604 ( .A(DW6[23]), .Y(n3717) );
    zmux21lb U1605 ( .A(n3716), .B(n3715), .S(n3324), .Y(UP_DW6[24]) );
    zivb U1606 ( .A(DW6[24]), .Y(n3715) );
    zmux21lb U1607 ( .A(n3714), .B(n3713), .S(n3941), .Y(UP_DW6[25]) );
    zivb U1608 ( .A(DW6[25]), .Y(n3713) );
    zmux21lb U1609 ( .A(n3712), .B(n3711), .S(n3324), .Y(UP_DW6[26]) );
    zivb U1610 ( .A(DW6[26]), .Y(n3711) );
    zmux21lb U1611 ( .A(n3710), .B(n3709), .S(n3941), .Y(UP_DW6[27]) );
    zivb U1612 ( .A(DW6[27]), .Y(n3709) );
    zmux21lb U1613 ( .A(n3708), .B(n3707), .S(n3324), .Y(UP_DW6[28]) );
    zivb U1614 ( .A(DW6[28]), .Y(n3707) );
    zmux21lb U1615 ( .A(n3706), .B(n3705), .S(n3941), .Y(UP_DW6[29]) );
    zivb U1616 ( .A(DW6[29]), .Y(n3705) );
    zmux21lb U1617 ( .A(n3704), .B(n3703), .S(n3941), .Y(UP_DW6[30]) );
    zivb U1618 ( .A(DW6[30]), .Y(n3703) );
    zivd U1619 ( .A(n3325), .Y(n3941) );
    zor2b U1620 ( .A(UP_LDW7), .B(QHSM[11]), .Y(n3325) );
    zmux21lb U1621 ( .A(n3099), .B(n3356), .S(n3537), .Y(UP_DW6[31]) );
    zivb U1622 ( .A(DW6[31]), .Y(n3356) );
    zan2b U1623 ( .A(INACT_COND), .B(n3324), .Y(n3537) );
    zivb U1624 ( .A(n3493), .Y(INACT_COND) );
    zivd U1625 ( .A(n3325), .Y(n3324) );
    zan3b U1626 ( .A(n3122), .B(n3118), .C(n3123), .Y(QHPARSING) );
    zivb U1627 ( .A(PHASENXT_idle), .Y(n3118) );
    zivb U1628 ( .A(n3649), .Y(n3086) );
    znd2b U1629 ( .A(n3906), .B(n3090), .Y(n3123) );
    zivb U1630 ( .A(n3122), .Y(QHSMNXT_13) );
    zivb U1631 ( .A(n3123), .Y(QHSMNXT_12) );
    zdffrb MULT_reg_1 ( .CK(PCICLK), .D(MULT588_1), .R(TRST_), .Q(MULT_1), 
        .QN(n3029) );
    zdffqrb MULT_reg_0 ( .CK(PCICLK), .D(MULT588_0), .R(TRST_), .Q(MULT_0) );
    zivb U1632 ( .A(MULT_0), .Y(MULT572_0) );
    zdffqrb TOTALBYTES_reg_14 ( .CK(PCICLK), .D(TOTALBYTES792_14), .R(TRST_), 
        .Q(TOTALBYTES_14) );
    zivb U1633 ( .A(TOTALBYTES_14), .Y(n3704) );
    zdffqrb TOTALBYTES_reg_13 ( .CK(PCICLK), .D(TOTALBYTES792_13), .R(TRST_), 
        .Q(TOTALBYTES_13) );
    zivb U1634 ( .A(TOTALBYTES_13), .Y(n3706) );
    zdffqrb TOTALBYTES_reg_12 ( .CK(PCICLK), .D(TOTALBYTES792_12), .R(TRST_), 
        .Q(TOTALBYTES_12) );
    zivb U1635 ( .A(TOTALBYTES_12), .Y(n3708) );
    zdffqrb TOTALBYTES_reg_11 ( .CK(PCICLK), .D(TOTALBYTES792_11), .R(TRST_), 
        .Q(TOTALBYTES_11) );
    zivb U1636 ( .A(TOTALBYTES_11), .Y(n3710) );
    zdffqrb TOTALBYTES_reg_10 ( .CK(PCICLK), .D(TOTALBYTES792_10), .R(TRST_), 
        .Q(TOTALBYTES_10) );
    zivb U1637 ( .A(TOTALBYTES_10), .Y(n3712) );
    zdffqrb TOTALBYTES_reg_9 ( .CK(PCICLK), .D(TOTALBYTES792_9), .R(TRST_), 
        .Q(TOTALBYTES_9) );
    zivb U1638 ( .A(TOTALBYTES_9), .Y(n3714) );
    zdffqrb TOTALBYTES_reg_8 ( .CK(PCICLK), .D(TOTALBYTES792_8), .R(TRST_), 
        .Q(TOTALBYTES_8) );
    zivb U1639 ( .A(TOTALBYTES_8), .Y(n3716) );
    zdffqrb TOTALBYTES_reg_7 ( .CK(PCICLK), .D(TOTALBYTES792_7), .R(TRST_), 
        .Q(TOTALBYTES_7) );
    zivb U1640 ( .A(TOTALBYTES_7), .Y(n3718) );
    zdffqrb TOTALBYTES_reg_6 ( .CK(PCICLK), .D(TOTALBYTES792_6), .R(TRST_), 
        .Q(TOTALBYTES_6) );
    zivb U1641 ( .A(TOTALBYTES_6), .Y(n3720) );
    zdffqrb TOTALBYTES_reg_5 ( .CK(PCICLK), .D(TOTALBYTES792_5), .R(TRST_), 
        .Q(TOTALBYTES_5) );
    zivb U1642 ( .A(TOTALBYTES_5), .Y(n3722) );
    zdffqrb TOTALBYTES_reg_4 ( .CK(PCICLK), .D(TOTALBYTES792_4), .R(TRST_), 
        .Q(TOTALBYTES_4) );
    zivb U1643 ( .A(TOTALBYTES_4), .Y(n3724) );
    zdffqrb TOTALBYTES_reg_3 ( .CK(PCICLK), .D(TOTALBYTES792_3), .R(TRST_), 
        .Q(TOTALBYTES_3) );
    zivb U1644 ( .A(TOTALBYTES_3), .Y(n3727) );
    zdffqrb TOTALBYTES_reg_2 ( .CK(PCICLK), .D(TOTALBYTES792_2), .R(TRST_), 
        .Q(TOTALBYTES_2) );
    zivb U1645 ( .A(TOTALBYTES_2), .Y(n3729) );
    zdffqrb TOTALBYTES_reg_1 ( .CK(PCICLK), .D(TOTALBYTES792_1), .R(TRST_), 
        .Q(TOTALBYTES_1) );
    zivb U1646 ( .A(TOTALBYTES_1), .Y(n3731) );
    zdffqrb TOTALBYTES_reg_0 ( .CK(PCICLK), .D(TOTALBYTES792_0), .R(TRST_), 
        .Q(TOTALBYTES_0) );
    zivb U1647 ( .A(TOTALBYTES_0), .Y(n3733) );
    zdffqb SBYTES_reg_6 ( .CK(PCICLK), .D(SBYTES962_6), .Q(UP_DW9[11]) );
    zdffqb SBYTES_reg_5 ( .CK(PCICLK), .D(SBYTES962_5), .Q(UP_DW9[10]) );
    zdffqb SBYTES_reg_4 ( .CK(PCICLK), .D(SBYTES962_4), .Q(UP_DW9[9]) );
    zdffqb SBYTES_reg_3 ( .CK(PCICLK), .D(SBYTES962_3), .Q(UP_DW9[8]) );
    zdffqb SBYTES_reg_2 ( .CK(PCICLK), .D(SBYTES962_2), .Q(UP_DW9[7]) );
    zdffqb SBYTES_reg_1 ( .CK(PCICLK), .D(SBYTES962_1), .Q(UP_DW9[6]) );
    zdffqb SBYTES_reg_0 ( .CK(PCICLK), .D(SBYTES962_0), .Q(UP_DW9[5]) );
    zdffqb CPAGE_reg_2 ( .CK(PCICLK), .D(CPAGE1173_2), .Q(CPAGE_2) );
    zivb U1648 ( .A(CPAGE_2), .Y(n3735) );
    zdffqb CPAGE_reg_1 ( .CK(PCICLK), .D(CPAGE1173_1), .Q(CPAGE_1) );
    zivb U1649 ( .A(CPAGE_1), .Y(n3737) );
    zdffqb CPROGMASK_reg_7 ( .CK(PCICLK), .D(CPROGMASK1402_7), .Q(UP_DW8[7])
         );
    zivb U1650 ( .A(UP_DW8[7]), .Y(n3668) );
    zdffqb CPROGMASK_reg_6 ( .CK(PCICLK), .D(CPROGMASK1402_6), .Q(UP_DW8[6])
         );
    zivb U1651 ( .A(UP_DW8[6]), .Y(n3664) );
    zdffqb CPROGMASK_reg_5 ( .CK(PCICLK), .D(CPROGMASK1402_5), .Q(UP_DW8[5])
         );
    zivb U1652 ( .A(UP_DW8[5]), .Y(n3669) );
    zdffqb CPROGMASK_reg_4 ( .CK(PCICLK), .D(CPROGMASK1402_4), .Q(UP_DW8[4])
         );
    zivb U1653 ( .A(UP_DW8[4]), .Y(n3665) );
    zdffqb CPROGMASK_reg_3 ( .CK(PCICLK), .D(CPROGMASK1402_3), .Q(UP_DW8[3])
         );
    zivb U1654 ( .A(UP_DW8[3]), .Y(n3666) );
    zdffqb CPROGMASK_reg_2 ( .CK(PCICLK), .D(CPROGMASK1402_2), .Q(UP_DW8[2])
         );
    zivb U1655 ( .A(UP_DW8[2]), .Y(n3670) );
    zdffqb CPROGMASK_reg_1 ( .CK(PCICLK), .D(CPROGMASK1402_1), .Q(UP_DW8[1])
         );
    zivb U1656 ( .A(UP_DW8[1]), .Y(n3667) );
    zdffqb CPROGMASK_reg_0 ( .CK(PCICLK), .D(CPROGMASK1402_0), .Q(UP_DW8[0])
         );
    zivb U1657 ( .A(UP_DW8[0]), .Y(n3526) );
    zdffqb FRAMETAG_reg_4 ( .CK(PCICLK), .D(FRAMETAG1470_4), .Q(UP_DW9[4]) );
    zdffqb FRAMETAG_reg_3 ( .CK(PCICLK), .D(FRAMETAG1470_3), .Q(UP_DW9[3]) );
    zdffqb FRAMETAG_reg_2 ( .CK(PCICLK), .D(FRAMETAG1470_2), .Q(UP_DW9[2]) );
    zdffqb FRAMETAG_reg_1 ( .CK(PCICLK), .D(FRAMETAG1470_1), .Q(UP_DW9[1]) );
    zdffqb FRAMETAG_reg_0 ( .CK(PCICLK), .D(FRAMETAG1470_0), .Q(UP_DW9[0]) );
    zdffb CURQTDPTR_reg_31 ( .CK(PCICLK), .D(CURQTDPTR1736_31), .Q(UP_DW3[31]), 
        .QN(n3142) );
    zdffb CURQTDPTR_reg_30 ( .CK(PCICLK), .D(CURQTDPTR1736_30), .Q(UP_DW3[30]), 
        .QN(n3148) );
    zdffb CURQTDPTR_reg_29 ( .CK(PCICLK), .D(CURQTDPTR1736_29), .Q(UP_DW3[29]), 
        .QN(n3152) );
    zdffb CURQTDPTR_reg_28 ( .CK(PCICLK), .D(CURQTDPTR1736_28), .Q(UP_DW3[28]), 
        .QN(n3156) );
    zdffb CURQTDPTR_reg_27 ( .CK(PCICLK), .D(CURQTDPTR1736_27), .Q(UP_DW3[27]), 
        .QN(n3160) );
    zdffb CURQTDPTR_reg_26 ( .CK(PCICLK), .D(CURQTDPTR1736_26), .Q(UP_DW3[26]), 
        .QN(n3164) );
    zdffb CURQTDPTR_reg_25 ( .CK(PCICLK), .D(CURQTDPTR1736_25), .Q(UP_DW3[25]), 
        .QN(n3168) );
    zdffb CURQTDPTR_reg_24 ( .CK(PCICLK), .D(CURQTDPTR1736_24), .Q(UP_DW3[24]), 
        .QN(n3172) );
    zdffb CURQTDPTR_reg_23 ( .CK(PCICLK), .D(CURQTDPTR1736_23), .Q(UP_DW3[23]), 
        .QN(n3176) );
    zdffb CURQTDPTR_reg_22 ( .CK(PCICLK), .D(CURQTDPTR1736_22), .Q(UP_DW3[22]), 
        .QN(n3180) );
    zdffb CURQTDPTR_reg_21 ( .CK(PCICLK), .D(CURQTDPTR1736_21), .Q(UP_DW3[21]), 
        .QN(n3184) );
    zdffb CURQTDPTR_reg_20 ( .CK(PCICLK), .D(CURQTDPTR1736_20), .Q(UP_DW3[20]), 
        .QN(n3188) );
    zdffb CURQTDPTR_reg_19 ( .CK(PCICLK), .D(CURQTDPTR1736_19), .Q(UP_DW3[19]), 
        .QN(n3192) );
    zdffb CURQTDPTR_reg_18 ( .CK(PCICLK), .D(CURQTDPTR1736_18), .Q(UP_DW3[18]), 
        .QN(n3196) );
    zdffb CURQTDPTR_reg_17 ( .CK(PCICLK), .D(CURQTDPTR1736_17), .Q(UP_DW3[17]), 
        .QN(n3200) );
    zdffb CURQTDPTR_reg_16 ( .CK(PCICLK), .D(CURQTDPTR1736_16), .Q(UP_DW3[16]), 
        .QN(n3204) );
    zdffb CURQTDPTR_reg_15 ( .CK(PCICLK), .D(CURQTDPTR1736_15), .Q(UP_DW3[15]), 
        .QN(n3208) );
    zdffb CURQTDPTR_reg_14 ( .CK(PCICLK), .D(CURQTDPTR1736_14), .Q(UP_DW3[14]), 
        .QN(n3212) );
    zdffb CURQTDPTR_reg_13 ( .CK(PCICLK), .D(CURQTDPTR1736_13), .Q(UP_DW3[13]), 
        .QN(n3216) );
    zdffb CURQTDPTR_reg_12 ( .CK(PCICLK), .D(CURQTDPTR1736_12), .Q(UP_DW3[12]), 
        .QN(n3220) );
    zdffb CURQTDPTR_reg_11 ( .CK(PCICLK), .D(CURQTDPTR1736_11), .Q(UP_DW3[11]), 
        .QN(n3224) );
    zdffb CURQTDPTR_reg_10 ( .CK(PCICLK), .D(CURQTDPTR1736_10), .Q(UP_DW3[10]), 
        .QN(n3228) );
    zdffb CURQTDPTR_reg_9 ( .CK(PCICLK), .D(CURQTDPTR1736_9), .Q(UP_DW3[9]), 
        .QN(n3232) );
    zdffb CURQTDPTR_reg_8 ( .CK(PCICLK), .D(CURQTDPTR1736_8), .Q(UP_DW3[8]), 
        .QN(n3236) );
    zdffb CURQTDPTR_reg_7 ( .CK(PCICLK), .D(CURQTDPTR1736_7), .Q(UP_DW3[7]), 
        .QN(n3240) );
    zdffb CURQTDPTR_reg_6 ( .CK(PCICLK), .D(CURQTDPTR1736_6), .Q(UP_DW3[6]), 
        .QN(n3244) );
    zdffb CURQTDPTR_reg_5 ( .CK(PCICLK), .D(CURQTDPTR1736_5), .Q(UP_DW3[5]), 
        .QN(n3248) );
    zdffqb OVERWBOFFSET_reg_11 ( .CK(PCICLK), .D(OVERWBOFFSET2136_11), .Q(
        UP_DW7[11]) );
    zdffqb OVERWBOFFSET_reg_10 ( .CK(PCICLK), .D(OVERWBOFFSET2136_10), .Q(
        UP_DW7[10]) );
    zdffqb OVERWBOFFSET_reg_9 ( .CK(PCICLK), .D(OVERWBOFFSET2136_9), .Q(UP_DW7
        [9]) );
    zdffqb OVERWBOFFSET_reg_8 ( .CK(PCICLK), .D(OVERWBOFFSET2136_8), .Q(UP_DW7
        [8]) );
    zdffqb OVERWBOFFSET_reg_7 ( .CK(PCICLK), .D(OVERWBOFFSET2136_7), .Q(UP_DW7
        [7]) );
    zdffqb OVERWBOFFSET_reg_6 ( .CK(PCICLK), .D(OVERWBOFFSET2136_6), .Q(UP_DW7
        [6]) );
    zdffqb OVERWBOFFSET_reg_5 ( .CK(PCICLK), .D(OVERWBOFFSET2136_5), .Q(UP_DW7
        [5]) );
    zdffqb OVERWBOFFSET_reg_4 ( .CK(PCICLK), .D(OVERWBOFFSET2136_4), .Q(UP_DW7
        [4]) );
    zdffqb OVERWBOFFSET_reg_3 ( .CK(PCICLK), .D(OVERWBOFFSET2136_3), .Q(UP_DW7
        [3]) );
    zdffqb OVERWBOFFSET_reg_2 ( .CK(PCICLK), .D(OVERWBOFFSET2136_2), .Q(UP_DW7
        [2]) );
    zdffqb OVERWBOFFSET_reg_1 ( .CK(PCICLK), .D(OVERWBOFFSET2136_1), .Q(UP_DW7
        [1]) );
    zdffqb OVERWBOFFSET_reg_0 ( .CK(PCICLK), .D(OVERWBOFFSET2136_0), .Q(UP_DW7
        [0]) );
    zivb U1658 ( .A(QHSM[9]), .Y(n3689) );
    zdffqrb HCI_PRESOF_T_reg ( .CK(PCICLK), .D(HCI_PRESOF_T1608), .R(TRST_), 
        .Q(HCI_PRESOF_T) );
    zdffqrb QHSM_reg_13 ( .CK(PCICLK), .D(QHSMNXT_13), .R(TRST_), .Q(QHSM[13])
         );
    zivb U1659 ( .A(QHSM[13]), .Y(n3783) );
    zivc U1660 ( .A(QHSM[0]), .Y(n3127) );
    zdffqrb PARSEQHEND_reg ( .CK(PCICLK), .D(PARSEQHEND_PRE), .R(TRST_), .Q(
        PARSEQHEND) );
    zdffqrb QEOT_reg ( .CK(PCICLK), .D(QEOT2302), .R(TRST_), .Q(QEOT) );
    zdffqrb_ UP_CACHE1_reg ( .CK(PCICLK), .D(QHSM[2]), .R(TRST_), .Q(UP_CACHE1
        ) );
    zivb U1661 ( .A(UP_CACHE1), .Y(n3702) );
    zivc U1662 ( .A(TRAN_CMD[14]), .Y(n3104) );
    zdffqrb QHSM_reg_7 ( .CK(PCICLK), .D(QHSMNXT_7), .R(TRST_), .Q(QHSM[7]) );
    zivb U1663 ( .A(QHSM[7]), .Y(n3654) );
    zdffqb ACTIVE_reg ( .CK(PCICLK), .D(ACTIVE_NXT), .Q(ACTIVE) );
    zivb U1664 ( .A(ACTIVE), .Y(n3590) );
    zdffqrb QHSM_reg_6 ( .CK(PCICLK), .D(PHASENXT_outcyc), .R(TRST_), .Q(QHSM
        [6]) );
    zivb U1665 ( .A(QHSM[6]), .Y(n3690) );
    zdffqrb QHSM_reg_8 ( .CK(PCICLK), .D(QHSMNXT_8), .R(TRST_), .Q(QHSM[8]) );
    zivb U1666 ( .A(QHSM[8]), .Y(n3775) );
    zdffrb PING_ERR_reg ( .CK(PCICLK), .D(PING_ERR1014), .R(TRST_), .Q(
        PING_ERR), .QN(n3829) );
    zdffqrb IMMEDRETRY_reg ( .CK(PCICLK), .D(IMMEDRETRY1571), .R(TRST_), .Q(
        IMMEDRETRY) );
    zivb U1667 ( .A(IMMEDRETRY), .Y(n3491) );
    zdffqrb QHSM_reg_1 ( .CK(PCICLK), .D(QHSMNXT_1), .R(TRST_), .Q(QHSM[1]) );
    zivb U1668 ( .A(QHSM[1]), .Y(n3596) );
    zdffqrb_ QRXERR_CUR_reg ( .CK(PCICLK), .D(QRXERR_CUR1646), .R(TRST_), .Q(
        QRXERR) );
    zdffb XACTERR_reg ( .CK(PCICLK), .D(XACTERR1308), .QN(n3535) );
    zdffqrb_ UP_CACHE2_reg ( .CK(PCICLK), .D(QHSM[11]), .R(TRST_), .Q(UP_LDW7)
         );
    zdffqrb QHSM_reg_10 ( .CK(PCICLK), .D(QHSMNXT_10), .R(TRST_), .Q(QHSM[10])
         );
    zivb U1669 ( .A(QHSM[10]), .Y(n3093) );
    zdffqrb CACHE_INVALID_reg ( .CK(PCICLK), .D(CACHE_INVALID1964), .R(TRST_), 
        .Q(CACHE_INVALID) );
    zdffqrb QHSM_reg_3 ( .CK(PCICLK), .D(QHSMNXT_3), .R(TRST_), .Q(QHSM[3]) );
    zivb U1670 ( .A(QHSM[3]), .Y(n3600) );
    zdffrb CACHE_MODIFY_reg ( .CK(PCICLK), .D(CACHE_MODIFY502), .R(TRST_), .Q(
        CACHE_MODIFY), .QN(n3588) );
    zdffb MISUF_reg ( .CK(PCICLK), .D(MISUF1318), .QN(n3601) );
    zdffqrb QHIOCINT_T_reg ( .CK(EHCIFLOW_PCLK), .D(QHIOCINT_T2339), .R(TRST_), 
        .Q(QHIOCINT_T) );
    zivb U1671 ( .A(QHIOCINT_T), .Y(n3135) );
    zdffqrb QHSM_reg_4 ( .CK(PCICLK), .D(QHSMNXT_4), .R(TRST_), .Q(QHSM[4]) );
    zivb U1672 ( .A(QHSM[4]), .Y(n3777) );
    zdffqrb QHSM_reg_5 ( .CK(PCICLK), .D(QHSMNXT_5), .R(TRST_), .Q(QHSM[5]) );
    zivb U1673 ( .A(QHSM[5]), .Y(n3595) );
    zdffqrb QCMDSTART_EOT_reg ( .CK(PCICLK), .D(QCMDSTART_EOT2265), .R(TRST_), 
        .Q(QCMDSTART_EOT) );
    zivb U1674 ( .A(QCMDSTART_EOT), .Y(n3102) );
    zdffrb SPLITXSTATE_OLD_reg ( .CK(PCICLK), .D(SPLITXSTATE_OLD1378), .R(
        TRST_), .QN(n3764) );
    zdffrb LENGTMAX_reg ( .CK(PCICLK), .D(LENGTMAX867), .R(TRST_), .QN(n3641)
         );
    zdffqrb QHERRINT_reg ( .CK(EHCIFLOW_PCLK), .D(QHERRINT2450), .R(TRST_), 
        .Q(QHERRINT) );
    zdffqrb QHIOCINT_reg ( .CK(EHCIFLOW_PCLK), .D(QHIOCINT2376), .R(TRST_), 
        .Q(QHIOCINT) );
    zdffqrb QHSM_reg_11 ( .CK(PCICLK), .D(PHASENXT_resultwb), .R(TRST_), .Q(
        QHSM[11]) );
    zivb U1675 ( .A(QHSM[11]), .Y(n3640) );
    zdffqrb QHERRINT_T_reg ( .CK(EHCIFLOW_PCLK), .D(QHERRINT_T2413), .R(TRST_), 
        .Q(QHERRINT_T) );
    zivb U1676 ( .A(QHERRINT_T), .Y(n3320) );
    zdffqb QTDHALT_reg ( .CK(PCICLK), .D(n2908), .Q(QTDHALT) );
    zivb U1677 ( .A(QTDHALT), .Y(n3827) );
    zdffb DT_reg ( .CK(PCICLK), .D(DT1086), .Q(DT), .QN(n3099) );
    zivb U1678 ( .A(QHSM[2]), .Y(n3652) );
    znr2b U1679 ( .A(INACT_COND), .B(n3702), .Y(UP_LDW3) );
    zdffb CERR_reg_1 ( .CK(PCICLK), .D(CERR1251_1), .Q(CERR_1), .QN(n3085) );
    znr3d U1680 ( .A(RECOVERYMODE), .B(n3633), .C(n2889), .Y(n2868) );
    znr5b U1681 ( .A(n2891), .B(n3538), .C(n2921), .D(n3743), .E(n3633), .Y(
        n2869) );
    znr2b U1682 ( .A(n3642), .B(n3598), .Y(n2870) );
    znr2d U1683 ( .A(n3769), .B(n2927), .Y(n2871) );
    znr2d U1684 ( .A(n3810), .B(n2927), .Y(n2872) );
    znr4b U1685 ( .A(QHSM[7]), .B(n3595), .C(n3532), .D(n3653), .Y(n2873) );
    znr4b U1686 ( .A(QHSM[8]), .B(n3690), .C(n3106), .D(n3653), .Y(n2874) );
    znr4b U1687 ( .A(QHSM[5]), .B(n3654), .C(n3532), .D(n3653), .Y(n2875) );
    znr3d U1688 ( .A(n2930), .B(n3783), .C(n3781), .Y(n2876) );
    znr2b U1689 ( .A(UP_DW6[8]), .B(n3125), .Y(TRAN_CMD[7]) );
    zan2b U1690 ( .A(TOTAL_SBYTES_10), .B(n3329), .Y(n2878) );
    zan2b U1691 ( .A(TOTAL_SBYTES_1), .B(n3329), .Y(n2879) );
    zan2b U1692 ( .A(TOTAL_SBYTES_0), .B(n3329), .Y(n2880) );
    znr3b U1693 ( .A(n3786), .B(n3751), .C(n3753), .Y(n2881) );
    znr2d U1694 ( .A(GEN_PERR), .B(n3105), .Y(n2882) );
    znr2d U1695 ( .A(n3602), .B(n3807), .Y(n2883) );
    znr3b U1696 ( .A(n3778), .B(n3124), .C(n2926), .Y(n2884) );
    znr2b U1697 ( .A(n2927), .B(n3818), .Y(n2885) );
    znr2b U1698 ( .A(n3817), .B(n2927), .Y(n2886) );
    znr6b U1699 ( .A(n3590), .B(n3641), .C(n3642), .D(BABBLE), .E(SPD), .F(
        QRXERR), .Y(n2887) );
    zoa21b U1700 ( .A(n3100), .B(n3648), .C(RECOVERYMODE), .Y(n2888) );
    znr2d U1701 ( .A(n3845), .B(n3846), .Y(n2889) );
    zan8b U1702 ( .A(n3691), .B(n3692), .C(n3693), .D(n3694), .E(n3695), .F(
        n3696), .G(n3697), .H(n3698), .Y(n2890) );
    znr3b U1703 ( .A(CPAGE_0), .B(CPAGE_1), .C(n3735), .Y(n2891) );
    znr2b U1704 ( .A(RXDATA0), .B(RXDATA1), .Y(n2892) );
    znr2b U1705 ( .A(CERR_1), .B(CERR_0), .Y(n2893) );
    zaoi21b U1706 ( .A(RXNYET), .B(n2890), .C(RXPIDERR), .Y(n2894) );
    zaoi21b U1707 ( .A(RXACK), .B(n3023), .C(RXNAK), .Y(n2895) );
    znr2b U1708 ( .A(n3814), .B(n3785), .Y(n2896) );
    zmux21hb U1709 ( .A(n2878), .B(DW1[26]), .S(n2923), .Y(MAXLEN[10]) );
    zmux21hb U1710 ( .A(TOTALBYTES_REAL_9), .B(DW1[25]), .S(n2923), .Y(MAXLEN
        [9]) );
    zmux21hb U1711 ( .A(TOTALBYTES_REAL_8), .B(DW1[24]), .S(n2923), .Y(MAXLEN
        [8]) );
    zmux21hb U1712 ( .A(TOTALBYTES_REAL_7), .B(DW1[23]), .S(n2923), .Y(MAXLEN
        [7]) );
    zmux21hb U1713 ( .A(TOTALBYTES_REAL_6), .B(DW1[22]), .S(n2923), .Y(MAXLEN
        [6]) );
    zmux21hb U1714 ( .A(TOTALBYTES_REAL_5), .B(DW1[21]), .S(n2923), .Y(MAXLEN
        [5]) );
    zmux21hb U1715 ( .A(TOTALBYTES_REAL_4), .B(DW1[20]), .S(n2923), .Y(MAXLEN
        [4]) );
    zmux21hb U1716 ( .A(TOTALBYTES_REAL_3), .B(DW1[19]), .S(n2923), .Y(MAXLEN
        [3]) );
    zmux21hb U1717 ( .A(TOTALBYTES_REAL_2), .B(DW1[18]), .S(n2923), .Y(MAXLEN
        [2]) );
    zmux21hb U1718 ( .A(n2879), .B(DW1[17]), .S(n2923), .Y(MAXLEN[1]) );
    zmux21hb U1719 ( .A(n2880), .B(DW1[16]), .S(LENGTMAX_PRE), .Y(MAXLEN[0])
         );
    zmux21hb U1720 ( .A(n3832), .B(DW6[6]), .S(LDPARM), .Y(n2908) );
    zdffqb CPAGE_reg_0 ( .CK(PCICLK), .D(CPAGE1173_0), .Q(CPAGE_0) );
    zivb U1721 ( .A(CPAGE_0), .Y(n3739) );
    zdffqb CERR_reg_0 ( .CK(PCICLK), .D(CERR1251_0), .Q(CERR_0) );
    zivb U1722 ( .A(CERR_0), .Y(n3828) );
    zmux21lb U1723 ( .A(TRAN_CMD[42]), .B(ACTLEN[2]), .S(n2519), .Y(n2909) );
    zmux21lb U1724 ( .A(TRAN_CMD[40]), .B(ACTLEN[0]), .S(n2519), .Y(n2910) );
    zmux21lb U1725 ( .A(TRAN_CMD[41]), .B(ACTLEN[1]), .S(n2519), .Y(n2911) );
    znd2b U1726 ( .A(DW9[9]), .B(n3358), .Y(n2912) );
    znd2b U1727 ( .A(DW9[8]), .B(n3358), .Y(n2913) );
    znd2b U1728 ( .A(DW9[10]), .B(n3358), .Y(n2914) );
    znd2b U1729 ( .A(DW9[7]), .B(n3358), .Y(n2915) );
    znd2b U1730 ( .A(DW9[11]), .B(n3358), .Y(n2916) );
    znd2b U1731 ( .A(DW9[5]), .B(n3358), .Y(n2917) );
    znd2b U1732 ( .A(DW9[6]), .B(n3358), .Y(n2918) );
    zivb U1733 ( .A(n3917), .Y(TOTALBYTES_REAL_2) );
    znd2b U1734 ( .A(TOTAL_SBYTES_2), .B(n3329), .Y(n3917) );
    zivb U1735 ( .A(n3915), .Y(TOTALBYTES_REAL_4) );
    znd2b U1736 ( .A(TOTAL_SBYTES_4), .B(n3329), .Y(n3915) );
    zivb U1737 ( .A(n3916), .Y(TOTALBYTES_REAL_3) );
    znd2b U1738 ( .A(TOTAL_SBYTES_3), .B(n3329), .Y(n3916) );
    zivb U1739 ( .A(n3913), .Y(TOTALBYTES_REAL_6) );
    znd2b U1740 ( .A(TOTAL_SBYTES_6), .B(n3329), .Y(n3913) );
    zivb U1741 ( .A(n3914), .Y(TOTALBYTES_REAL_5) );
    znd2b U1742 ( .A(TOTAL_SBYTES_5), .B(n3329), .Y(n3914) );
    zivb U1743 ( .A(n3911), .Y(TOTALBYTES_REAL_8) );
    znd2b U1744 ( .A(TOTAL_SBYTES_8), .B(n3329), .Y(n3911) );
    zivb U1745 ( .A(n3912), .Y(TOTALBYTES_REAL_7) );
    znd2b U1746 ( .A(TOTAL_SBYTES_7), .B(n3329), .Y(n3912) );
    zivb U1747 ( .A(n3910), .Y(TOTALBYTES_REAL_9) );
    znd2b U1748 ( .A(TOTAL_SBYTES_9), .B(n3329), .Y(n3910) );
    znr2b U1749 ( .A(sub_451_carry_14), .B(TOTALBYTES_14), .Y(n2919) );
    znr2b U1750 ( .A(sub_457_carry_14), .B(TOTALBYTES_REAL_14), .Y(n2920) );
    zivc U1751 ( .A(n3023), .Y(TRAN_CMD[9]) );
    ziv11b U1752 ( .A(n3023), .Y(UP_DW6[8]), .Z(n2921) );
    zor2b U1753 ( .A(n3063), .B(n3061), .Y(n2922) );
    znd2d U1754 ( .A(n3084), .B(n2922), .Y(n2923) );
    zivb U1755 ( .A(n2923), .Y(n3839) );
    znd2b U1756 ( .A(n3084), .B(n2922), .Y(LENGTMAX_PRE) );
    zoai2x4b U1757 ( .A(n3195), .B(n3927), .C(n3928), .D(n3196), .E(n3197), 
        .F(n3930), .G(n3198), .H(n3932), .Y(CURQTDPTR1736_18) );
    zoai2x4b U1758 ( .A(n3239), .B(n3927), .C(n3141), .D(n3240), .E(n3241), 
        .F(n3929), .G(n3242), .H(n3932), .Y(CURQTDPTR1736_7) );
    zoai2x4b U1759 ( .A(n3183), .B(n3927), .C(n3928), .D(n3184), .E(n3185), 
        .F(n3930), .G(n3186), .H(n3932), .Y(CURQTDPTR1736_21) );
    zoai2x4b U1760 ( .A(n3219), .B(n3927), .C(n3928), .D(n3220), .E(n3221), 
        .F(n3930), .G(n3222), .H(n3932), .Y(CURQTDPTR1736_12) );
    zoai2x4b U1761 ( .A(n3167), .B(n3927), .C(n3141), .D(n3168), .E(n3169), 
        .F(n3929), .G(n3170), .H(n3931), .Y(CURQTDPTR1736_25) );
    zoai2x4b U1762 ( .A(n3231), .B(n3927), .C(n3141), .D(n3232), .E(n3233), 
        .F(n3930), .G(n3234), .H(n3931), .Y(CURQTDPTR1736_9) );
    zor3d U1763 ( .A(n3133), .B(n3127), .C(n3815), .Y(n3927) );
    zoai2x4b U1764 ( .A(n3199), .B(n3140), .C(n3141), .D(n3200), .E(n3201), 
        .F(n3144), .G(n3202), .H(n3146), .Y(CURQTDPTR1736_17) );
    zoai2x4b U1765 ( .A(n3151), .B(n3140), .C(n3141), .D(n3152), .E(n3153), 
        .F(n3144), .G(n3154), .H(n3146), .Y(CURQTDPTR1736_29) );
    zoai2x4b U1766 ( .A(n3211), .B(n3140), .C(n3928), .D(n3212), .E(n3213), 
        .F(n3144), .G(n3214), .H(n3146), .Y(CURQTDPTR1736_14) );
    zoai2x4b U1767 ( .A(n3175), .B(n3140), .C(n3928), .D(n3176), .E(n3177), 
        .F(n3144), .G(n3178), .H(n3146), .Y(CURQTDPTR1736_23) );
    zoai2x4b U1768 ( .A(n3223), .B(n3140), .C(n3141), .D(n3224), .E(n3225), 
        .F(n3144), .G(n3226), .H(n3146), .Y(CURQTDPTR1736_11) );
    zoai2x4b U1769 ( .A(n3163), .B(n3140), .C(n3928), .D(n3164), .E(n3165), 
        .F(n3144), .G(n3166), .H(n3146), .Y(CURQTDPTR1736_26) );
    zor3d U1770 ( .A(n3133), .B(n3127), .C(n3815), .Y(n3140) );
    zor3d U1771 ( .A(n3133), .B(n3127), .C(n3815), .Y(n3926) );
    zivb U1772 ( .A(n3813), .Y(n3815) );
    zivb U1773 ( .A(n3793), .Y(n2924) );
    zivd U1774 ( .A(DWCNT[1]), .Y(n3793) );
    zivb U1775 ( .A(n3799), .Y(n2925) );
    zivd U1776 ( .A(DWCNT[2]), .Y(n3799) );
    zivb U1777 ( .A(n3090), .Y(n2926) );
    zor2b U1778 ( .A(n2926), .B(n3834), .Y(n3122) );
    zor2b U1779 ( .A(GEN_PERR), .B(n3569), .Y(n3811) );
    zivb U1780 ( .A(GEN_PERR), .Y(n3090) );
    zor2b U1781 ( .A(GEN_PERR), .B(n3521), .Y(n3115) );
    zor2b U1782 ( .A(GEN_PERR), .B(n3495), .Y(n3114) );
    zao21b U1783 ( .A(n3779), .B(n3780), .C(GEN_PERR), .Y(n3111) );
    zbfd U1784 ( .A(n3128), .Y(n2927) );
    zbfb U1785 ( .A(n3128), .Y(n2928) );
    zor2b U1786 ( .A(n2927), .B(n3770), .Y(n3772) );
    zor2b U1787 ( .A(n3767), .B(n2927), .Y(n3807) );
    zivb U1788 ( .A(n2927), .Y(n3766) );
    zor2b U1789 ( .A(NXTISSTSWB), .B(n2928), .Y(n3597) );
    zor2b U1790 ( .A(n3753), .B(n2928), .Y(n3360) );
    zor2b U1791 ( .A(n3768), .B(QH_PARSE_GO), .Y(n3128) );
    zbfd U1792 ( .A(QHSM_12), .Y(QHSM[12]) );
    zbfd U1793 ( .A(QHSM_12), .Y(n2931) );
    zbfb U1794 ( .A(QHSM_12), .Y(n2930) );
    zivc U1795 ( .A(n2930), .Y(QHDWNUM[0]) );
    zdffqrb QHSM_reg_12 ( .CK(PCICLK), .D(QHSMNXT_12), .R(TRST_), .Q(QHSM_12)
         );
    zbfd U1796 ( .A(DW6[8]), .Y(n2932) );
    zan2b U1797 ( .A(UP_DW6[8]), .B(n3103), .Y(TRAN_CMD[1]) );
    zor2b U1798 ( .A(UP_DW6[8]), .B(n3126), .Y(TRAN_CMD[104]) );
    zaoi222b U1799 ( .A(OVERWBOFFSET_P2090_12), .B(n3608), .C(n3609), .D(
        CUROFFSET_T_12), .E(OVERWBOFFSET_P2070_12), .F(n2932), .Y(n3607) );
    zxo2b U1800 ( .A(TRAN_CMD[14]), .B(n2932), .Y(n3771) );
    zan3b U1801 ( .A(n2932), .B(QHSM[3]), .C(n3556), .Y(n3555) );
    zor2b U1802 ( .A(n2932), .B(n3100), .Y(n3805) );
    zor2b U1803 ( .A(n2932), .B(n2893), .Y(n3553) );
    znd3b U1804 ( .A(n2932), .B(RXMDATA), .C(n3358), .Y(n3548) );
    zor2b U1805 ( .A(TRAN_CMD[6]), .B(n2932), .Y(n3748) );
    zao21b U1806 ( .A(n2932), .B(TRAN_CMD[14]), .C(n3100), .Y(n2519) );
    zbfb U1807 ( .A(DW1[12]), .Y(TRAN_CMD[13]) );
    zbfb U1808 ( .A(DW2[23]), .Y(TRAN_CMD[15]) );
    zbfb U1809 ( .A(DW2[24]), .Y(TRAN_CMD[16]) );
    zbfb U1810 ( .A(DW2[25]), .Y(TRAN_CMD[17]) );
    zbfb U1811 ( .A(DW2[26]), .Y(TRAN_CMD[18]) );
    zbfb U1812 ( .A(DW2[27]), .Y(TRAN_CMD[19]) );
    zbfb U1813 ( .A(DW2[28]), .Y(TRAN_CMD[20]) );
    zbfb U1814 ( .A(DW2[29]), .Y(TRAN_CMD[21]) );
    zbfb U1815 ( .A(DW2[16]), .Y(TRAN_CMD[22]) );
    zbfb U1816 ( .A(DW2[17]), .Y(TRAN_CMD[23]) );
    zbfb U1817 ( .A(DW2[18]), .Y(TRAN_CMD[24]) );
    zbfb U1818 ( .A(DW2[19]), .Y(TRAN_CMD[25]) );
    zbfb U1819 ( .A(DW2[20]), .Y(TRAN_CMD[26]) );
    zbfb U1820 ( .A(DW2[21]), .Y(TRAN_CMD[27]) );
    zbfb U1821 ( .A(DW2[22]), .Y(TRAN_CMD[28]) );
    zbfb U1822 ( .A(DW1[8]), .Y(TRAN_CMD[29]) );
    zbfb U1823 ( .A(DW1[9]), .Y(TRAN_CMD[30]) );
    zbfb U1824 ( .A(DW1[10]), .Y(TRAN_CMD[31]) );
    zbfb U1825 ( .A(DW1[11]), .Y(TRAN_CMD[32]) );
    zbfb U1826 ( .A(DW1[0]), .Y(TRAN_CMD[33]) );
    zbfb U1827 ( .A(DW1[1]), .Y(TRAN_CMD[34]) );
    zbfb U1828 ( .A(DW1[2]), .Y(TRAN_CMD[35]) );
    zbfb U1829 ( .A(DW1[3]), .Y(TRAN_CMD[36]) );
    zbfb U1830 ( .A(DW1[4]), .Y(TRAN_CMD[37]) );
    zbfb U1831 ( .A(DW1[5]), .Y(TRAN_CMD[38]) );
    zbfb U1832 ( .A(DW1[6]), .Y(TRAN_CMD[39]) );
    zbfb U1833 ( .A(QHCIMWR), .Y(QHCIADR[3]) );
    zor2b U1834 ( .A(QHSM[13]), .B(n2930), .Y(QHCIMWR) );
    zbfb U1835 ( .A(QHDWNUM[2]), .Y(QHDWNUM[1]) );
    zivb U1836 ( .A(QHCIMWR), .Y(QHDWNUM[2]) );
    zbfb U1837 ( .A(QHDWNUM[3]), .Y(QHCIADR[2]) );
    zivb U1838 ( .A(n3797), .Y(QHDWNUM[3]) );
    zbfb U1839 ( .A(UP_LDW9), .Y(UP_LDW8) );
    zor2b U1840 ( .A(UP_LDW7), .B(UP_LDW3), .Y(UP_LDW9) );
    zbfb U1841 ( .A(DW9[12]), .Y(UP_DW9[12]) );
    zbfb U1842 ( .A(DW9[13]), .Y(UP_DW9[13]) );
    zbfb U1843 ( .A(DW9[14]), .Y(UP_DW9[14]) );
    zbfb U1844 ( .A(DW9[15]), .Y(UP_DW9[15]) );
    zbfb U1845 ( .A(DW9[16]), .Y(UP_DW9[16]) );
    zbfb U1846 ( .A(DW9[17]), .Y(UP_DW9[17]) );
    zbfb U1847 ( .A(DW9[18]), .Y(UP_DW9[18]) );
    zbfb U1848 ( .A(DW9[19]), .Y(UP_DW9[19]) );
    zbfb U1849 ( .A(DW9[20]), .Y(UP_DW9[20]) );
    zbfb U1850 ( .A(DW9[21]), .Y(UP_DW9[21]) );
    zbfb U1851 ( .A(DW9[22]), .Y(UP_DW9[22]) );
    zbfb U1852 ( .A(DW9[23]), .Y(UP_DW9[23]) );
    zbfb U1853 ( .A(DW9[24]), .Y(UP_DW9[24]) );
    zbfb U1854 ( .A(DW9[25]), .Y(UP_DW9[25]) );
    zbfb U1855 ( .A(DW9[26]), .Y(UP_DW9[26]) );
    zbfb U1856 ( .A(DW9[27]), .Y(UP_DW9[27]) );
    zbfb U1857 ( .A(DW9[28]), .Y(UP_DW9[28]) );
    zbfb U1858 ( .A(DW9[29]), .Y(UP_DW9[29]) );
    zbfb U1859 ( .A(DW9[30]), .Y(UP_DW9[30]) );
    zbfb U1860 ( .A(DW9[31]), .Y(UP_DW9[31]) );
    zbfb U1861 ( .A(DW8[12]), .Y(UP_DW8[12]) );
    zbfb U1862 ( .A(DW8[13]), .Y(UP_DW8[13]) );
    zbfb U1863 ( .A(DW8[14]), .Y(UP_DW8[14]) );
    zbfb U1864 ( .A(DW8[15]), .Y(UP_DW8[15]) );
    zbfb U1865 ( .A(DW8[16]), .Y(UP_DW8[16]) );
    zbfb U1866 ( .A(DW8[17]), .Y(UP_DW8[17]) );
    zbfb U1867 ( .A(DW8[18]), .Y(UP_DW8[18]) );
    zbfb U1868 ( .A(DW8[19]), .Y(UP_DW8[19]) );
    zbfb U1869 ( .A(DW8[20]), .Y(UP_DW8[20]) );
    zbfb U1870 ( .A(DW8[21]), .Y(UP_DW8[21]) );
    zbfb U1871 ( .A(DW8[22]), .Y(UP_DW8[22]) );
    zbfb U1872 ( .A(DW8[23]), .Y(UP_DW8[23]) );
    zbfb U1873 ( .A(DW8[24]), .Y(UP_DW8[24]) );
    zbfb U1874 ( .A(DW8[25]), .Y(UP_DW8[25]) );
    zbfb U1875 ( .A(DW8[26]), .Y(UP_DW8[26]) );
    zbfb U1876 ( .A(DW8[27]), .Y(UP_DW8[27]) );
    zbfb U1877 ( .A(DW8[28]), .Y(UP_DW8[28]) );
    zbfb U1878 ( .A(DW8[29]), .Y(UP_DW8[29]) );
    zbfb U1879 ( .A(DW8[30]), .Y(UP_DW8[30]) );
    zbfb U1880 ( .A(DW8[31]), .Y(UP_DW8[31]) );
    zbfb U1881 ( .A(DW7[12]), .Y(UP_DW7[12]) );
    zbfb U1882 ( .A(DW7[13]), .Y(UP_DW7[13]) );
    zbfb U1883 ( .A(DW7[14]), .Y(UP_DW7[14]) );
    zbfb U1884 ( .A(DW7[15]), .Y(UP_DW7[15]) );
    zbfb U1885 ( .A(DW7[16]), .Y(UP_DW7[16]) );
    zbfb U1886 ( .A(DW7[17]), .Y(UP_DW7[17]) );
    zbfb U1887 ( .A(DW7[18]), .Y(UP_DW7[18]) );
    zbfb U1888 ( .A(DW7[19]), .Y(UP_DW7[19]) );
    zbfb U1889 ( .A(DW7[20]), .Y(UP_DW7[20]) );
    zbfb U1890 ( .A(DW7[21]), .Y(UP_DW7[21]) );
    zbfb U1891 ( .A(DW7[22]), .Y(UP_DW7[22]) );
    zbfb U1892 ( .A(DW7[23]), .Y(UP_DW7[23]) );
    zbfb U1893 ( .A(DW7[24]), .Y(UP_DW7[24]) );
    zbfb U1894 ( .A(DW7[25]), .Y(UP_DW7[25]) );
    zbfb U1895 ( .A(DW7[26]), .Y(UP_DW7[26]) );
    zbfb U1896 ( .A(DW7[27]), .Y(UP_DW7[27]) );
    zbfb U1897 ( .A(DW7[28]), .Y(UP_DW7[28]) );
    zbfb U1898 ( .A(DW7[29]), .Y(UP_DW7[29]) );
    zbfb U1899 ( .A(DW7[30]), .Y(UP_DW7[30]) );
    zbfb U1900 ( .A(DW7[31]), .Y(UP_DW7[31]) );
    zivb U1901 ( .A(n2932), .Y(n3023) );
    zbfb U1902 ( .A(DW6[9]), .Y(UP_DW6[9]) );
    zbfb U1903 ( .A(DW6[15]), .Y(UP_DW6[15]) );
    zbfb U1904 ( .A(QHSM[0]), .Y(QHIDLE) );
    zan2b U1905 ( .A(UP_DW9[5]), .B(ACTLEN[0]), .Y(add_508_carry_1) );
    zxo2b U1906 ( .A(UP_DW9[5]), .B(ACTLEN[0]), .Y(SBYTES966_0) );
    zxo2b U1907 ( .A(add_919_carry_12), .B(CUROFFSET_T_12), .Y(
        OVERWBOFFSET_P2070_12) );
    zan2b U1908 ( .A(UP_DW7[11]), .B(add_922_carry_11), .Y(
        OVERWBOFFSET_P2090_12) );
    zxo2b U1909 ( .A(UP_DW7[11]), .B(add_922_carry_11), .Y(
        OVERWBOFFSET_P2090_11) );
    zan2b U1910 ( .A(TRAN_CMD[83]), .B(add_919_carry_11), .Y(add_919_carry_12)
         );
    zxo2b U1911 ( .A(TRAN_CMD[83]), .B(add_919_carry_11), .Y(
        OVERWBOFFSET_P2070_11) );
    zan2b U1912 ( .A(UP_DW7[11]), .B(r481_carry_11), .Y(CUROFFSET_T_12) );
    zxo2b U1913 ( .A(UP_DW7[11]), .B(r481_carry_11), .Y(TRAN_CMD[83]) );
    zan2b U1914 ( .A(UP_DW7[10]), .B(r481_carry_10), .Y(r481_carry_11) );
    zxo2b U1915 ( .A(UP_DW7[10]), .B(r481_carry_10), .Y(TRAN_CMD[82]) );
    zan2b U1916 ( .A(UP_DW7[9]), .B(r481_carry_9), .Y(r481_carry_10) );
    zxo2b U1917 ( .A(UP_DW7[9]), .B(r481_carry_9), .Y(TRAN_CMD[81]) );
    zan2b U1918 ( .A(UP_DW7[8]), .B(r481_carry_8), .Y(r481_carry_9) );
    zxo2b U1919 ( .A(UP_DW7[8]), .B(r481_carry_8), .Y(TRAN_CMD[80]) );
    zan2b U1920 ( .A(UP_DW7[7]), .B(r481_carry_7), .Y(r481_carry_8) );
    zxo2b U1921 ( .A(UP_DW7[7]), .B(r481_carry_7), .Y(TRAN_CMD[79]) );
    zan2b U1922 ( .A(UP_DW7[0]), .B(MAXLEN[0]), .Y(add_922_carry_1) );
    zxo2b U1923 ( .A(UP_DW7[0]), .B(MAXLEN[0]), .Y(OVERWBOFFSET_P2090_0) );
    zan2b U1924 ( .A(TRAN_CMD[72]), .B(ACTLEN[0]), .Y(add_919_carry_1) );
    zxo2b U1925 ( .A(TRAN_CMD[72]), .B(ACTLEN[0]), .Y(OVERWBOFFSET_P2070_0) );
    zan2b U1926 ( .A(UP_DW9[5]), .B(UP_DW7[0]), .Y(r481_carry_1) );
    zxo2b U1927 ( .A(UP_DW9[5]), .B(UP_DW7[0]), .Y(TRAN_CMD[72]) );
    zxn2b U1928 ( .A(sub_457_carry_14), .B(TOTALBYTES_REAL_14), .Y(
        VIR_TOTALBYTES_14) );
    zor2b U1929 ( .A(sub_457_carry_13), .B(TOTALBYTES_REAL_13), .Y(
        sub_457_carry_14) );
    zxn2b U1930 ( .A(sub_457_carry_13), .B(TOTALBYTES_REAL_13), .Y(
        VIR_TOTALBYTES_13) );
    zor2b U1931 ( .A(sub_457_carry_12), .B(TOTALBYTES_REAL_12), .Y(
        sub_457_carry_13) );
    zxn2b U1932 ( .A(sub_457_carry_12), .B(TOTALBYTES_REAL_12), .Y(
        VIR_TOTALBYTES_12) );
    zor2b U1933 ( .A(sub_457_carry_11), .B(TOTALBYTES_REAL_11), .Y(
        sub_457_carry_12) );
    zxn2b U1934 ( .A(sub_457_carry_11), .B(TOTALBYTES_REAL_11), .Y(
        VIR_TOTALBYTES_11) );
    zor2b U1935 ( .A(n2880), .B(n2910), .Y(sub_457_carry_1) );
    zxn2b U1936 ( .A(n2880), .B(n2910), .Y(VIR_TOTALBYTES_0) );
    zxn2b U1937 ( .A(sub_451_carry_14), .B(TOTALBYTES_14), .Y(TOTAL_SBYTES_14)
         );
    zor2b U1938 ( .A(sub_451_carry_13), .B(TOTALBYTES_13), .Y(sub_451_carry_14
        ) );
    zxn2b U1939 ( .A(sub_451_carry_13), .B(TOTALBYTES_13), .Y(TOTAL_SBYTES_13)
         );
    zor2b U1940 ( .A(sub_451_carry_12), .B(TOTALBYTES_12), .Y(sub_451_carry_13
        ) );
    zxn2b U1941 ( .A(sub_451_carry_12), .B(TOTALBYTES_12), .Y(TOTAL_SBYTES_12)
         );
    zor2b U1942 ( .A(sub_451_carry_11), .B(TOTALBYTES_11), .Y(sub_451_carry_12
        ) );
    zxn2b U1943 ( .A(sub_451_carry_11), .B(TOTALBYTES_11), .Y(TOTAL_SBYTES_11)
         );
    zor2b U1944 ( .A(sub_451_carry_10), .B(TOTALBYTES_10), .Y(sub_451_carry_11
        ) );
    zxn2b U1945 ( .A(sub_451_carry_10), .B(TOTALBYTES_10), .Y(TOTAL_SBYTES_10)
         );
    zor2b U1946 ( .A(sub_451_carry_9), .B(TOTALBYTES_9), .Y(sub_451_carry_10)
         );
    zxn2b U1947 ( .A(sub_451_carry_9), .B(TOTALBYTES_9), .Y(TOTAL_SBYTES_9) );
    zor2b U1948 ( .A(sub_451_carry_8), .B(TOTALBYTES_8), .Y(sub_451_carry_9)
         );
    zxn2b U1949 ( .A(sub_451_carry_8), .B(TOTALBYTES_8), .Y(TOTAL_SBYTES_8) );
    zor2b U1950 ( .A(sub_451_carry_7), .B(TOTALBYTES_7), .Y(sub_451_carry_8)
         );
    zxn2b U1951 ( .A(sub_451_carry_7), .B(TOTALBYTES_7), .Y(TOTAL_SBYTES_7) );
    zor2b U1952 ( .A(TOTALBYTES_0), .B(n2917), .Y(sub_451_carry_1) );
    zxn2b U1953 ( .A(TOTALBYTES_0), .B(n2917), .Y(TOTAL_SBYTES_0) );
    zymx24hb U1954 ( .A1(TRAN_CMD[46]), .A2(TRAN_CMD[45]), .A3(TRAN_CMD[44]), 
        .A4(TRAN_CMD[43]), .B1(ACTLEN[6]), .B2(ACTLEN[5]), .B3(ACTLEN[4]), 
        .B4(ACTLEN[3]), .S(n2519), .Y1(MINUEND_6), .Y2(MINUEND_5), .Y3(
        MINUEND_4), .Y4(MINUEND_3) );
    zymx24hb U1955 ( .A1(TRAN_CMD[50]), .A2(TRAN_CMD[49]), .A3(TRAN_CMD[48]), 
        .A4(TRAN_CMD[47]), .B1(ACTLEN[10]), .B2(ACTLEN[9]), .B3(ACTLEN[8]), 
        .B4(ACTLEN[7]), .S(n2519), .Y1(MINUEND_10), .Y2(MINUEND_9), .Y3(
        MINUEND_8), .Y4(MINUEND_7) );
    zdffqsd QHSM_reg_0 ( .CK(PCICLK), .D(PHASENXT_idle), .S(TRST_), .Q(QHSM[0]
        ) );
    zdffqrd SPLITXSTATE_reg ( .CK(PCICLK), .D(SPLITXSTATE1341), .R(TRST_), .Q(
        TRAN_CMD[14]) );
    zdffqrd QHSM_reg_2 ( .CK(PCICLK), .D(QHSMNXT_2), .R(TRST_), .Q(QHSM[2]) );
    znd2d U1956 ( .A(TOTALBYTES_REAL_2), .B(n3056), .Y(n3050) );
    znr3d U1957 ( .A(n3032), .B(TOTALBYTES_REAL_14), .C(TOTALBYTES_REAL_13), 
        .Y(n3084) );
    znd2d U1958 ( .A(n3050), .B(n3049), .Y(n3078) );
    znr2d U1959 ( .A(n3077), .B(n3074), .Y(n3075) );
    znr2d U1960 ( .A(n3079), .B(n3076), .Y(n3077) );
    znr2d U1961 ( .A(n3081), .B(n3078), .Y(n3079) );
    znr2d U1962 ( .A(n2879), .B(n3082), .Y(n3083) );
    zfa1b add_922_U1_5 ( .A(MAXLEN[5]), .B(UP_DW7[5]), .CI(add_922_carry_5), 
        .CO(add_922_carry_6), .S(OVERWBOFFSET_P2090_5) );
    zfa1b add_922_U1_4 ( .A(MAXLEN[4]), .B(UP_DW7[4]), .CI(add_922_carry_4), 
        .CO(add_922_carry_5), .S(OVERWBOFFSET_P2090_4) );
    zfa1b add_922_U1_3 ( .A(MAXLEN[3]), .B(UP_DW7[3]), .CI(add_922_carry_3), 
        .CO(add_922_carry_4), .S(OVERWBOFFSET_P2090_3) );
    zfa1b add_922_U1_10 ( .A(MAXLEN[10]), .B(UP_DW7[10]), .CI(add_922_carry_10
        ), .CO(add_922_carry_11), .S(OVERWBOFFSET_P2090_10) );
    zfa1b add_922_U1_9 ( .A(MAXLEN[9]), .B(UP_DW7[9]), .CI(add_922_carry_9), 
        .CO(add_922_carry_10), .S(OVERWBOFFSET_P2090_9) );
    zfa1b add_922_U1_2 ( .A(MAXLEN[2]), .B(UP_DW7[2]), .CI(add_922_carry_2), 
        .CO(add_922_carry_3), .S(OVERWBOFFSET_P2090_2) );
    zfa1b add_922_U1_7 ( .A(MAXLEN[7]), .B(UP_DW7[7]), .CI(add_922_carry_7), 
        .CO(add_922_carry_8), .S(OVERWBOFFSET_P2090_7) );
    zfa1b add_922_U1_8 ( .A(MAXLEN[8]), .B(UP_DW7[8]), .CI(add_922_carry_8), 
        .CO(add_922_carry_9), .S(OVERWBOFFSET_P2090_8) );
    zfa1b add_922_U1_6 ( .A(MAXLEN[6]), .B(UP_DW7[6]), .CI(add_922_carry_6), 
        .CO(add_922_carry_7), .S(OVERWBOFFSET_P2090_6) );
    zfa1b add_922_U1_1 ( .A(MAXLEN[1]), .B(UP_DW7[1]), .CI(add_922_carry_1), 
        .CO(add_922_carry_2), .S(OVERWBOFFSET_P2090_1) );
    zfa1b sub_451_U2_6 ( .A(TOTALBYTES_6), .B(n2916), .CI(sub_451_carry_6), 
        .CO(sub_451_carry_7), .S(TOTAL_SBYTES_6) );
    zfa1b sub_451_U2_1 ( .A(TOTALBYTES_1), .B(n2918), .CI(sub_451_carry_1), 
        .CO(sub_451_carry_2), .S(TOTAL_SBYTES_1) );
    zfa1b sub_451_U2_5 ( .A(TOTALBYTES_5), .B(n2914), .CI(sub_451_carry_5), 
        .CO(sub_451_carry_6), .S(TOTAL_SBYTES_5) );
    zfa1b sub_451_U2_3 ( .A(TOTALBYTES_3), .B(n2913), .CI(sub_451_carry_3), 
        .CO(sub_451_carry_4), .S(TOTAL_SBYTES_3) );
    zfa1b sub_451_U2_2 ( .A(TOTALBYTES_2), .B(n2915), .CI(sub_451_carry_2), 
        .CO(sub_451_carry_3), .S(TOTAL_SBYTES_2) );
    zfa1b sub_451_U2_4 ( .A(TOTALBYTES_4), .B(n2912), .CI(sub_451_carry_4), 
        .CO(sub_451_carry_5), .S(TOTAL_SBYTES_4) );
    zfa1b sub_457_U2_6 ( .A(TOTALBYTES_REAL_6), .B(sub_457_B_not_6), .CI(
        sub_457_carry_6), .CO(sub_457_carry_7), .S(VIR_TOTALBYTES_6) );
    zfa1b sub_457_U2_8 ( .A(TOTALBYTES_REAL_8), .B(sub_457_B_not_8), .CI(
        sub_457_carry_8), .CO(sub_457_carry_9), .S(VIR_TOTALBYTES_8) );
    zfa1b sub_457_U2_10 ( .A(n2878), .B(sub_457_B_not_10), .CI(
        sub_457_carry_10), .CO(sub_457_carry_11), .S(VIR_TOTALBYTES_10) );
    zfa1b sub_457_U2_9 ( .A(TOTALBYTES_REAL_9), .B(sub_457_B_not_9), .CI(
        sub_457_carry_9), .CO(sub_457_carry_10), .S(VIR_TOTALBYTES_9) );
    zfa1b sub_457_U2_1 ( .A(n2879), .B(n2911), .CI(sub_457_carry_1), .CO(
        sub_457_carry_2), .S(VIR_TOTALBYTES_1) );
    zfa1b sub_457_U2_7 ( .A(TOTALBYTES_REAL_7), .B(sub_457_B_not_7), .CI(
        sub_457_carry_7), .CO(sub_457_carry_8), .S(VIR_TOTALBYTES_7) );
    zfa1b sub_457_U2_5 ( .A(TOTALBYTES_REAL_5), .B(sub_457_B_not_5), .CI(
        sub_457_carry_5), .CO(sub_457_carry_6), .S(VIR_TOTALBYTES_5) );
    zfa1b sub_457_U2_3 ( .A(TOTALBYTES_REAL_3), .B(sub_457_B_not_3), .CI(
        sub_457_carry_3), .CO(sub_457_carry_4), .S(VIR_TOTALBYTES_3) );
    zfa1b sub_457_U2_2 ( .A(TOTALBYTES_REAL_2), .B(n2909), .CI(sub_457_carry_2
        ), .CO(sub_457_carry_3), .S(VIR_TOTALBYTES_2) );
    zfa1b sub_457_U2_4 ( .A(TOTALBYTES_REAL_4), .B(sub_457_B_not_4), .CI(
        sub_457_carry_4), .CO(sub_457_carry_5), .S(VIR_TOTALBYTES_4) );
    zfa1b add_508_U1_5 ( .A(ACTLEN[5]), .B(UP_DW9[10]), .CI(add_508_carry_5), 
        .CO(add_508_carry_6), .S(SBYTES966_5) );
    zfa1b add_508_U1_4 ( .A(ACTLEN[4]), .B(UP_DW9[9]), .CI(add_508_carry_4), 
        .CO(add_508_carry_5), .S(SBYTES966_4) );
    zfa1b add_508_U1_3 ( .A(ACTLEN[3]), .B(UP_DW9[8]), .CI(add_508_carry_3), 
        .CO(add_508_carry_4), .S(SBYTES966_3) );
    zfa1b add_508_U1_2 ( .A(ACTLEN[2]), .B(UP_DW9[7]), .CI(add_508_carry_2), 
        .CO(add_508_carry_3), .S(SBYTES966_2) );
    zfa1b add_508_U1_1 ( .A(ACTLEN[1]), .B(UP_DW9[6]), .CI(add_508_carry_1), 
        .CO(add_508_carry_2), .S(SBYTES966_1) );
    zfa1b add_919_U1_5 ( .A(ACTLEN[5]), .B(TRAN_CMD[77]), .CI(add_919_carry_5), 
        .CO(add_919_carry_6), .S(OVERWBOFFSET_P2070_5) );
    zfa1b add_919_U1_4 ( .A(ACTLEN[4]), .B(TRAN_CMD[76]), .CI(add_919_carry_4), 
        .CO(add_919_carry_5), .S(OVERWBOFFSET_P2070_4) );
    zfa1b add_919_U1_3 ( .A(ACTLEN[3]), .B(TRAN_CMD[75]), .CI(add_919_carry_3), 
        .CO(add_919_carry_4), .S(OVERWBOFFSET_P2070_3) );
    zfa1b add_919_U1_10 ( .A(ACTLEN[10]), .B(TRAN_CMD[82]), .CI(
        add_919_carry_10), .CO(add_919_carry_11), .S(OVERWBOFFSET_P2070_10) );
    zfa1b add_919_U1_9 ( .A(ACTLEN[9]), .B(TRAN_CMD[81]), .CI(add_919_carry_9), 
        .CO(add_919_carry_10), .S(OVERWBOFFSET_P2070_9) );
    zfa1b add_919_U1_2 ( .A(ACTLEN[2]), .B(TRAN_CMD[74]), .CI(add_919_carry_2), 
        .CO(add_919_carry_3), .S(OVERWBOFFSET_P2070_2) );
    zfa1b add_919_U1_7 ( .A(ACTLEN[7]), .B(TRAN_CMD[79]), .CI(add_919_carry_7), 
        .CO(add_919_carry_8), .S(OVERWBOFFSET_P2070_7) );
    zfa1b add_919_U1_8 ( .A(ACTLEN[8]), .B(TRAN_CMD[80]), .CI(add_919_carry_8), 
        .CO(add_919_carry_9), .S(OVERWBOFFSET_P2070_8) );
    zfa1b add_919_U1_6 ( .A(ACTLEN[6]), .B(TRAN_CMD[78]), .CI(add_919_carry_6), 
        .CO(add_919_carry_7), .S(OVERWBOFFSET_P2070_6) );
    zfa1b add_919_U1_1 ( .A(ACTLEN[1]), .B(TRAN_CMD[73]), .CI(add_919_carry_1), 
        .CO(add_919_carry_2), .S(OVERWBOFFSET_P2070_1) );
    zfa1b r481_U1_5 ( .A(UP_DW7[5]), .B(UP_DW9[10]), .CI(r481_carry_5), .CO(
        r481_carry_6), .S(TRAN_CMD[77]) );
    zfa1b r481_U1_4 ( .A(UP_DW7[4]), .B(UP_DW9[9]), .CI(r481_carry_4), .CO(
        r481_carry_5), .S(TRAN_CMD[76]) );
    zfa1b r481_U1_3 ( .A(UP_DW7[3]), .B(UP_DW9[8]), .CI(r481_carry_3), .CO(
        r481_carry_4), .S(TRAN_CMD[75]) );
    zfa1b r481_U1_2 ( .A(UP_DW7[2]), .B(UP_DW9[7]), .CI(r481_carry_2), .CO(
        r481_carry_3), .S(TRAN_CMD[74]) );
    zfa1b r481_U1_6 ( .A(UP_DW7[6]), .B(UP_DW9[11]), .CI(r481_carry_6), .CO(
        r481_carry_7), .S(TRAN_CMD[78]) );
    zfa1b r481_U1_1 ( .A(UP_DW7[1]), .B(UP_DW9[6]), .CI(r481_carry_1), .CO(
        r481_carry_2), .S(TRAN_CMD[73]) );
    zao211b U1963 ( .A(n3086), .B(n3087), .C(n3088), .D(n3089), .Y(
        PHASENXT_idle) );
    zind2d U1964 ( .A(DW1[12]), .B(DW1[13]), .Y(TRAN_CMD[6]) );
    zao211b U1965 ( .A(n3105), .B(n3106), .C(QHSM[9]), .D(n3107), .Y(QEOT2302)
         );
    zoai22d U1966 ( .A(n3116), .B(n3117), .C(n3118), .D(n3119), .Y(
        CACHE_INVALID1964) );
    zoa21d U1967 ( .A(QCMDSTART_EOT), .B(QCMDSTART), .C(n3124), .Y(
        QCMDSTART_EOT2265) );
    zao222b U1968 ( .A(DW6[14]), .B(n2927), .C(n2886), .D(CPAGE_2), .E(n2885), 
        .F(CPAGE1177_2), .Y(CPAGE1173_2) );
    zao222b U1969 ( .A(DW6[13]), .B(n2927), .C(n2886), .D(CPAGE_1), .E(n2885), 
        .F(CPAGE1177_1), .Y(CPAGE1173_1) );
    zao222b U1970 ( .A(DW6[12]), .B(n2927), .C(n2886), .D(CPAGE_0), .E(n2885), 
        .F(n3739), .Y(CPAGE1173_0) );
    zan4b U1971 ( .A(n3095), .B(n3127), .C(n3129), .D(n3130), .Y(
        QRXERR_CUR1646) );
    zao211b U1972 ( .A(DW6[0]), .B(n3934), .C(n3253), .D(n3254), .Y(QHCIADD[0]
        ) );
    zao211b U1973 ( .A(DW6[1]), .B(n3252), .C(n3255), .D(n3256), .Y(QHCIADD[1]
        ) );
    zao211b U1974 ( .A(DW6[2]), .B(n3933), .C(n3257), .D(n3258), .Y(QHCIADD[2]
        ) );
    zao211b U1975 ( .A(DW6[3]), .B(n3934), .C(n3259), .D(n3260), .Y(QHCIADD[3]
        ) );
    zao211b U1976 ( .A(DW6[4]), .B(n3252), .C(n3261), .D(n3262), .Y(QHCIADD[4]
        ) );
    zao211b U1977 ( .A(DW6[5]), .B(n3252), .C(n3263), .D(n3264), .Y(QHCIADD[5]
        ) );
    zao211b U1978 ( .A(DW6[6]), .B(n3933), .C(n3265), .D(n3266), .Y(QHCIADD[6]
        ) );
    zao211b U1979 ( .A(DW6[7]), .B(n3934), .C(n3267), .D(n3268), .Y(QHCIADD[7]
        ) );
    zao211b U1980 ( .A(TRAN_CMD[9]), .B(n3252), .C(n3269), .D(n3270), .Y(
        QHCIADD[8]) );
    zao211b U1981 ( .A(DW6[9]), .B(n3933), .C(n3271), .D(n3272), .Y(QHCIADD[9]
        ) );
    zao211b U1982 ( .A(DW6[10]), .B(n3934), .C(n3273), .D(n3274), .Y(QHCIADD
        [10]) );
    zao211b U1983 ( .A(DW6[11]), .B(n3933), .C(n3275), .D(n3276), .Y(QHCIADD
        [11]) );
    zao211b U1984 ( .A(DW6[12]), .B(n3934), .C(n3277), .D(n3278), .Y(QHCIADD
        [12]) );
    zao211b U1985 ( .A(DW6[13]), .B(n3252), .C(n3279), .D(n3280), .Y(QHCIADD
        [13]) );
    zao211b U1986 ( .A(DW6[14]), .B(n3933), .C(n3281), .D(n3282), .Y(QHCIADD
        [14]) );
    zao211b U1987 ( .A(DW6[15]), .B(n3934), .C(n3283), .D(n3284), .Y(QHCIADD
        [15]) );
    zao211b U1988 ( .A(DW6[16]), .B(n3252), .C(n3285), .D(n3286), .Y(QHCIADD
        [16]) );
    zao211b U1989 ( .A(DW6[17]), .B(n3933), .C(n3287), .D(n3288), .Y(QHCIADD
        [17]) );
    zao211b U1990 ( .A(DW6[18]), .B(n3934), .C(n3289), .D(n3290), .Y(QHCIADD
        [18]) );
    zao211b U1991 ( .A(DW6[19]), .B(n3252), .C(n3291), .D(n3292), .Y(QHCIADD
        [19]) );
    zao211b U1992 ( .A(DW6[20]), .B(n3252), .C(n3293), .D(n3294), .Y(QHCIADD
        [20]) );
    zao211b U1993 ( .A(DW6[21]), .B(n3933), .C(n3295), .D(n3296), .Y(QHCIADD
        [21]) );
    zao211b U1994 ( .A(DW6[22]), .B(n3934), .C(n3297), .D(n3298), .Y(QHCIADD
        [22]) );
    zao211b U1995 ( .A(DW6[23]), .B(n3933), .C(n3299), .D(n3300), .Y(QHCIADD
        [23]) );
    zao211b U1996 ( .A(DW6[24]), .B(n3934), .C(n3301), .D(n3302), .Y(QHCIADD
        [24]) );
    zao211b U1997 ( .A(DW6[25]), .B(n3252), .C(n3303), .D(n3304), .Y(QHCIADD
        [25]) );
    zao211b U1998 ( .A(DW6[26]), .B(n3933), .C(n3305), .D(n3306), .Y(QHCIADD
        [26]) );
    zao211b U1999 ( .A(DW6[27]), .B(n3934), .C(n3307), .D(n3308), .Y(QHCIADD
        [27]) );
    zao211b U2000 ( .A(DW6[28]), .B(n3252), .C(n3309), .D(n3310), .Y(QHCIADD
        [28]) );
    zao211b U2001 ( .A(DW6[29]), .B(n3252), .C(n3311), .D(n3312), .Y(QHCIADD
        [29]) );
    zao211b U2002 ( .A(DW6[30]), .B(n3933), .C(n3313), .D(n3314), .Y(QHCIADD
        [30]) );
    zao211b U2003 ( .A(DW6[31]), .B(n3934), .C(n3315), .D(n3316), .Y(QHCIADD
        [31]) );
    zao222b U2004 ( .A(n2871), .B(UP_DW9[11]), .C(n3322), .D(DW9[11]), .E(
        n3323), .F(SBYTES966_6), .Y(SBYTES962_6) );
    zao222b U2005 ( .A(UP_DW9[10]), .B(n2871), .C(n3322), .D(DW9[10]), .E(
        SBYTES966_5), .F(n3323), .Y(SBYTES962_5) );
    zao222b U2006 ( .A(UP_DW9[9]), .B(n2871), .C(n3322), .D(DW9[9]), .E(
        SBYTES966_4), .F(n3323), .Y(SBYTES962_4) );
    zao222b U2007 ( .A(UP_DW9[8]), .B(n2871), .C(n3322), .D(DW9[8]), .E(
        SBYTES966_3), .F(n3323), .Y(SBYTES962_3) );
    zao222b U2008 ( .A(UP_DW9[7]), .B(n2871), .C(n3322), .D(DW9[7]), .E(
        SBYTES966_2), .F(n3323), .Y(SBYTES962_2) );
    zao222b U2009 ( .A(UP_DW9[6]), .B(n2871), .C(n3322), .D(DW9[6]), .E(
        SBYTES966_1), .F(n3323), .Y(SBYTES962_1) );
    zao222b U2010 ( .A(UP_DW9[5]), .B(n2871), .C(n3322), .D(DW9[5]), .E(
        SBYTES966_0), .F(n3323), .Y(SBYTES962_0) );
    zao222b U2011 ( .A(n3326), .B(TOTALBYTES_14), .C(DW6[30]), .D(LDPARM), .E(
        VIR_TOTALBYTES_14), .F(n3328), .Y(TOTALBYTES792_14) );
    zao222b U2012 ( .A(n3326), .B(TOTALBYTES_13), .C(DW6[29]), .D(n3327), .E(
        VIR_TOTALBYTES_13), .F(n3328), .Y(TOTALBYTES792_13) );
    zao222b U2013 ( .A(n3326), .B(TOTALBYTES_12), .C(DW6[28]), .D(LDPARM), .E(
        VIR_TOTALBYTES_12), .F(n3328), .Y(TOTALBYTES792_12) );
    zao222b U2014 ( .A(n3326), .B(TOTALBYTES_11), .C(DW6[27]), .D(n3327), .E(
        VIR_TOTALBYTES_11), .F(n3328), .Y(TOTALBYTES792_11) );
    zao222b U2015 ( .A(n3326), .B(TOTALBYTES_10), .C(DW6[26]), .D(LDPARM), .E(
        VIR_TOTALBYTES_10), .F(n3328), .Y(TOTALBYTES792_10) );
    zao222b U2016 ( .A(n3326), .B(TOTALBYTES_9), .C(DW6[25]), .D(n3327), .E(
        VIR_TOTALBYTES_9), .F(n3328), .Y(TOTALBYTES792_9) );
    zao222b U2017 ( .A(n3326), .B(TOTALBYTES_8), .C(DW6[24]), .D(LDPARM), .E(
        VIR_TOTALBYTES_8), .F(n3328), .Y(TOTALBYTES792_8) );
    zao222b U2018 ( .A(n3326), .B(TOTALBYTES_7), .C(DW6[23]), .D(n3327), .E(
        VIR_TOTALBYTES_7), .F(n3328), .Y(TOTALBYTES792_7) );
    zao222b U2019 ( .A(n3326), .B(TOTALBYTES_6), .C(DW6[22]), .D(LDPARM), .E(
        VIR_TOTALBYTES_6), .F(n3328), .Y(TOTALBYTES792_6) );
    zao222b U2020 ( .A(n3326), .B(TOTALBYTES_5), .C(DW6[21]), .D(n3327), .E(
        VIR_TOTALBYTES_5), .F(n3328), .Y(TOTALBYTES792_5) );
    zao222b U2021 ( .A(n3326), .B(TOTALBYTES_4), .C(DW6[20]), .D(LDPARM), .E(
        VIR_TOTALBYTES_4), .F(n3328), .Y(TOTALBYTES792_4) );
    zao222b U2022 ( .A(n3326), .B(TOTALBYTES_3), .C(DW6[19]), .D(n3327), .E(
        VIR_TOTALBYTES_3), .F(n3328), .Y(TOTALBYTES792_3) );
    zao222b U2023 ( .A(n3326), .B(TOTALBYTES_2), .C(DW6[18]), .D(LDPARM), .E(
        VIR_TOTALBYTES_2), .F(n3328), .Y(TOTALBYTES792_2) );
    zao222b U2024 ( .A(n3326), .B(TOTALBYTES_1), .C(DW6[17]), .D(n3327), .E(
        VIR_TOTALBYTES_1), .F(n3328), .Y(TOTALBYTES792_1) );
    zao222b U2025 ( .A(n3326), .B(TOTALBYTES_0), .C(DW6[16]), .D(LDPARM), .E(
        VIR_TOTALBYTES_0), .F(n3328), .Y(TOTALBYTES792_0) );
    zao222b U2026 ( .A(UP_DW7[0]), .B(n3330), .C(DW7[0]), .D(n3331), .E(n3332), 
        .F(n3333), .Y(OVERWBOFFSET2136_0) );
    zao222b U2027 ( .A(UP_DW7[1]), .B(n3330), .C(DW7[1]), .D(n3331), .E(n3332), 
        .F(n3334), .Y(OVERWBOFFSET2136_1) );
    zao222b U2028 ( .A(UP_DW7[2]), .B(n3330), .C(DW7[2]), .D(n3331), .E(n3332), 
        .F(n3335), .Y(OVERWBOFFSET2136_2) );
    zao222b U2029 ( .A(UP_DW7[3]), .B(n3330), .C(DW7[3]), .D(n3331), .E(n3332), 
        .F(n3336), .Y(OVERWBOFFSET2136_3) );
    zao222b U2030 ( .A(UP_DW7[4]), .B(n3330), .C(DW7[4]), .D(n3331), .E(n3332), 
        .F(n3337), .Y(OVERWBOFFSET2136_4) );
    zao222b U2031 ( .A(UP_DW7[5]), .B(n3330), .C(DW7[5]), .D(n3331), .E(n3332), 
        .F(n3338), .Y(OVERWBOFFSET2136_5) );
    zao222b U2032 ( .A(UP_DW7[6]), .B(n3330), .C(DW7[6]), .D(n3331), .E(n3332), 
        .F(n3339), .Y(OVERWBOFFSET2136_6) );
    zao222b U2033 ( .A(UP_DW7[7]), .B(n3330), .C(DW7[7]), .D(n3331), .E(n3332), 
        .F(n3340), .Y(OVERWBOFFSET2136_7) );
    zao222b U2034 ( .A(UP_DW7[8]), .B(n3330), .C(DW7[8]), .D(n3331), .E(n3332), 
        .F(n3341), .Y(OVERWBOFFSET2136_8) );
    zao222b U2035 ( .A(UP_DW7[9]), .B(n3330), .C(DW7[9]), .D(n3331), .E(n3332), 
        .F(n3342), .Y(OVERWBOFFSET2136_9) );
    zao222b U2036 ( .A(UP_DW7[10]), .B(n3330), .C(DW7[10]), .D(n3331), .E(
        n3332), .F(n3343), .Y(OVERWBOFFSET2136_10) );
    zao222b U2037 ( .A(UP_DW7[11]), .B(n3330), .C(DW7[11]), .D(n3331), .E(
        n3332), .F(n3344), .Y(OVERWBOFFSET2136_11) );
    zao222b U2038 ( .A(DW8[0]), .B(n2927), .C(n3345), .D(n3346), .E(UP_DW8[0]), 
        .F(n3347), .Y(CPROGMASK1402_0) );
    zao222b U2039 ( .A(DW8[1]), .B(n2928), .C(n3345), .D(n3348), .E(UP_DW8[1]), 
        .F(n3347), .Y(CPROGMASK1402_1) );
    zao222b U2040 ( .A(DW8[2]), .B(n2927), .C(n3345), .D(n3349), .E(UP_DW8[2]), 
        .F(n3347), .Y(CPROGMASK1402_2) );
    zao222b U2041 ( .A(DW8[3]), .B(n2928), .C(n3345), .D(n3350), .E(UP_DW8[3]), 
        .F(n3347), .Y(CPROGMASK1402_3) );
    zao222b U2042 ( .A(DW8[4]), .B(n2927), .C(n3345), .D(n3351), .E(UP_DW8[4]), 
        .F(n3347), .Y(CPROGMASK1402_4) );
    zao222b U2043 ( .A(DW8[5]), .B(n2927), .C(n3345), .D(n3352), .E(UP_DW8[5]), 
        .F(n3347), .Y(CPROGMASK1402_5) );
    zao222b U2044 ( .A(DW8[6]), .B(n2927), .C(n3345), .D(n3353), .E(UP_DW8[6]), 
        .F(n3347), .Y(CPROGMASK1402_6) );
    zao222b U2045 ( .A(DW8[7]), .B(n2927), .C(n3345), .D(n3354), .E(UP_DW8[7]), 
        .F(n3347), .Y(CPROGMASK1402_7) );
    zao211b U2046 ( .A(DW7[31]), .B(n3362), .C(n3363), .D(n3364), .Y(TRAN_CMD
        [103]) );
    zao211b U2047 ( .A(DW7[30]), .B(n3362), .C(n3365), .D(n3366), .Y(TRAN_CMD
        [102]) );
    zao211b U2048 ( .A(DW7[29]), .B(n3362), .C(n3367), .D(n3368), .Y(TRAN_CMD
        [101]) );
    zao211b U2049 ( .A(DW7[28]), .B(n3362), .C(n3369), .D(n3370), .Y(TRAN_CMD
        [100]) );
    zao211b U2050 ( .A(n3362), .B(DW7[27]), .C(n3371), .D(n3372), .Y(TRAN_CMD
        [99]) );
    zao211b U2051 ( .A(DW7[26]), .B(n3362), .C(n3373), .D(n3374), .Y(TRAN_CMD
        [98]) );
    zao211b U2052 ( .A(DW7[25]), .B(n3362), .C(n3375), .D(n3376), .Y(TRAN_CMD
        [97]) );
    zao211b U2053 ( .A(DW7[24]), .B(n3362), .C(n3377), .D(n3378), .Y(TRAN_CMD
        [96]) );
    zao211b U2054 ( .A(DW7[23]), .B(n3362), .C(n3379), .D(n3380), .Y(TRAN_CMD
        [95]) );
    zao211b U2055 ( .A(DW7[22]), .B(n3362), .C(n3381), .D(n3382), .Y(TRAN_CMD
        [94]) );
    zao211b U2056 ( .A(DW7[21]), .B(n3362), .C(n3383), .D(n3384), .Y(TRAN_CMD
        [93]) );
    zao211b U2057 ( .A(DW7[20]), .B(n3362), .C(n3385), .D(n3386), .Y(TRAN_CMD
        [92]) );
    zao211b U2058 ( .A(DW7[19]), .B(n3362), .C(n3387), .D(n3388), .Y(TRAN_CMD
        [91]) );
    zao211b U2059 ( .A(DW7[18]), .B(n3362), .C(n3389), .D(n3390), .Y(TRAN_CMD
        [90]) );
    zao211b U2060 ( .A(DW7[17]), .B(n3362), .C(n3391), .D(n3392), .Y(TRAN_CMD
        [89]) );
    zao211b U2061 ( .A(DW7[16]), .B(n3362), .C(n3393), .D(n3394), .Y(TRAN_CMD
        [88]) );
    zao211b U2062 ( .A(DW7[15]), .B(n3362), .C(n3395), .D(n3396), .Y(TRAN_CMD
        [87]) );
    zao211b U2063 ( .A(DW7[14]), .B(n3362), .C(n3397), .D(n3398), .Y(TRAN_CMD
        [86]) );
    zao211b U2064 ( .A(DW7[13]), .B(n3362), .C(n3399), .D(n3400), .Y(TRAN_CMD
        [85]) );
    zao211b U2065 ( .A(DW7[12]), .B(n3362), .C(n3401), .D(n3402), .Y(TRAN_CMD
        [84]) );
    zan4b U2066 ( .A(n3490), .B(n3491), .C(n2887), .D(n2882), .Y(n3097) );
    zoa21d U2067 ( .A(UP_DW8[6]), .B(n3500), .C(n3354), .Y(n3499) );
    zoa21d U2068 ( .A(UP_DW8[5]), .B(n3502), .C(n3353), .Y(n3501) );
    zoa21d U2069 ( .A(UP_DW8[4]), .B(n3504), .C(n3352), .Y(n3503) );
    zoa21d U2070 ( .A(UP_DW8[3]), .B(n3506), .C(n3351), .Y(n3505) );
    zoa21d U2071 ( .A(UP_DW8[2]), .B(n3508), .C(n3350), .Y(n3507) );
    zoa21d U2072 ( .A(UP_DW8[1]), .B(n3510), .C(n3349), .Y(n3509) );
    zoa21d U2073 ( .A(UP_DW8[0]), .B(n3512), .C(n3348), .Y(n3511) );
    zoa21d U2074 ( .A(UP_DW8[7]), .B(n3514), .C(n3346), .Y(n3513) );
    znr8d U2075 ( .A(n3499), .B(n3501), .C(n3503), .D(n3505), .E(n3507), .F(
        n3509), .G(n3511), .H(n3513), .Y(n3515) );
    zoa21d U2076 ( .A(n3517), .B(n3518), .C(n3519), .Y(n3516) );
    zoa21d U2077 ( .A(n3522), .B(n3523), .C(n3524), .Y(n3521) );
    zoa21d U2078 ( .A(QHSM[6]), .B(QHSM[9]), .C(PHASENXT_resultwb), .Y(n3094)
         );
    zan2d U2079 ( .A(n2890), .B(n3103), .Y(n3528) );
    zoa21d U2080 ( .A(n3528), .B(n3530), .C(RXNYET), .Y(n3529) );
    zan4b U2081 ( .A(QH_ACT), .B(n3532), .C(EHCI_MAC_EOT), .D(n3533), .Y(n3531
        ) );
    zan4b U2082 ( .A(n3539), .B(n3540), .C(n3541), .D(n3542), .Y(n3538) );
    zan4b U2083 ( .A(n3545), .B(n3546), .C(n3547), .D(n3548), .Y(n3544) );
    zoa21d U2084 ( .A(n2892), .B(n2921), .C(n2895), .Y(n3549) );
    zan4b U2085 ( .A(IMMEDRETRY), .B(n3105), .C(n3553), .D(n3554), .Y(n3552)
         );
    zoa21d U2086 ( .A(n2889), .B(n3126), .C(n3558), .Y(n3557) );
    zoa21d U2087 ( .A(n3562), .B(n3563), .C(n3564), .Y(n3561) );
    zoa21d U2088 ( .A(IMMEDRETRY), .B(n2887), .C(n3566), .Y(n3565) );
    zoa21d U2089 ( .A(QHCIMWR), .B(n3573), .C(QHSM[10]), .Y(n3572) );
    zoa21d U2090 ( .A(ACTIVE), .B(INACT_COND), .C(n3575), .Y(n3574) );
    zoa21d U2091 ( .A(n2896), .B(n3577), .C(n3578), .Y(n3576) );
    zoa21d U2092 ( .A(QHSM[0]), .B(n3586), .C(QHSM[3]), .Y(n3585) );
    zoa21d U2093 ( .A(n3579), .B(n3587), .C(n3588), .Y(n3089) );
    zan4b U2094 ( .A(n3590), .B(QHSM[13]), .C(DW6[15]), .D(n3122), .Y(n3589)
         );
    zoa21d U2095 ( .A(PARSEQHEND), .B(n3133), .C(n3596), .Y(n3120) );
    zoa21d U2096 ( .A(n3522), .B(n3600), .C(n3601), .Y(n3599) );
    zoa21d U2097 ( .A(n3104), .B(n3603), .C(n3604), .Y(n3602) );
    zoa21d U2098 ( .A(n3605), .B(n3606), .C(n3133), .Y(n3355) );
    zoa21d U2099 ( .A(n2895), .B(n3104), .C(TRAN_CMD[6]), .Y(n3610) );
    zan4b U2100 ( .A(n3126), .B(ACTIVE), .C(n2894), .D(n3624), .Y(n3623) );
    zan4b U2101 ( .A(n2932), .B(n3626), .C(n3627), .D(n3100), .Y(n3625) );
    zor2d U2102 ( .A(n3631), .B(n3104), .Y(n3633) );
    zor5b U2103 ( .A(QHSM[3]), .B(QHSM[4]), .C(QHSM[0]), .D(n3638), .E(QHCIREQ
        ), .Y(n3639) );
    zor5b U2104 ( .A(QHSM[10]), .B(QHSM[9]), .C(QHSM[2]), .D(n3640), .E(n3639), 
        .Y(n3643) );
    zor3b U2105 ( .A(QHSM[10]), .B(n3573), .C(QHCIMWR), .Y(n3645) );
    zor3b U2106 ( .A(QHSM[2]), .B(QHSM[3]), .C(n3646), .Y(n3647) );
    zor3b U2107 ( .A(n3586), .B(n3127), .C(n3647), .Y(n3649) );
    zor3b U2108 ( .A(n3133), .B(n3649), .C(n2888), .Y(n3650) );
    zor3b U2109 ( .A(QHSM[3]), .B(QHSM[0]), .C(n3586), .Y(n3651) );
    zor3b U2110 ( .A(QHSM[2]), .B(n3651), .C(n3645), .Y(n3653) );
    zor3b U2111 ( .A(n3655), .B(n3656), .C(n3657), .Y(n3603) );
    zor3b U2112 ( .A(FRNUM[0]), .B(n3656), .C(n3657), .Y(n3658) );
    zor3b U2113 ( .A(FRNUM[1]), .B(n3655), .C(n3657), .Y(n3659) );
    zor3b U2114 ( .A(FRNUM[1]), .B(FRNUM[0]), .C(n3657), .Y(n3660) );
    zor3b U2115 ( .A(FRNUM[2]), .B(n3655), .C(n3656), .Y(n3661) );
    zor3b U2116 ( .A(FRNUM[2]), .B(FRNUM[0]), .C(n3656), .Y(n3662) );
    zivh U2117 ( .A(DW2[10]), .Y(n3508) );
    zor3b U2118 ( .A(FRNUM[2]), .B(FRNUM[1]), .C(n3655), .Y(n3663) );
    zor3b U2119 ( .A(FRNUM[2]), .B(FRNUM[1]), .C(FRNUM[0]), .Y(n3527) );
    zivh U2120 ( .A(DW2[8]), .Y(n3512) );
    zor3b U2121 ( .A(n3671), .B(n3672), .C(n3515), .Y(n3517) );
    zor5b U2122 ( .A(n3673), .B(n3674), .C(n3675), .D(n3676), .E(n3677), .Y(
        n3518) );
    zoai21d U2123 ( .A(n3679), .B(n3680), .C(n3358), .Y(n3678) );
    zivh U2124 ( .A(DW2[6]), .Y(n3682) );
    zivh U2125 ( .A(DW2[5]), .Y(n3683) );
    zivh U2126 ( .A(DW2[4]), .Y(n3684) );
    zor5b U2127 ( .A(QHSM[2]), .B(QHSM[0]), .C(n3600), .D(n3586), .E(n3646), 
        .Y(n3523) );
    zor4b U2128 ( .A(QHSM[10]), .B(n3689), .C(CACHEPHASE), .D(n3639), .Y(n3496
        ) );
    zor4b U2129 ( .A(QHSM[9]), .B(n3093), .C(CACHEPHASE), .D(n3639), .Y(n3498)
         );
    zor3b U2130 ( .A(BABBLE), .B(QRXERR), .C(n3494), .Y(n3497) );
    zor3b U2131 ( .A(DW6[1]), .B(n3578), .C(n3644), .Y(n3493) );
    zor3b U2132 ( .A(n3628), .B(n3630), .C(n3948), .Y(n3744) );
    zor3b U2133 ( .A(n3746), .B(n3948), .C(n3628), .Y(n3407) );
    zor3b U2134 ( .A(n3747), .B(n3745), .C(n3630), .Y(n3405) );
    zor3b U2135 ( .A(n3746), .B(n3747), .C(n3745), .Y(n3403) );
    zor4b U2136 ( .A(BABBLE), .B(n3530), .C(n3544), .D(n3129), .Y(n3749) );
    zor3b U2137 ( .A(n3766), .B(n3648), .C(n3631), .Y(n3765) );
    zor3b U2138 ( .A(n3129), .B(n3771), .C(n3767), .Y(n3770) );
    zor3b U2139 ( .A(n2893), .B(n3774), .C(n3753), .Y(n3773) );
    zor4b U2140 ( .A(QHSM[6]), .B(n3775), .C(n3106), .D(n3653), .Y(n3776) );
    zor4b U2141 ( .A(QHSM[1]), .B(QHSM[0]), .C(n3777), .D(n3647), .Y(n3778) );
    zor4b U2142 ( .A(QHSM[4]), .B(QHSM[0]), .C(n3596), .D(n3647), .Y(n3571) );
    zor5b U2143 ( .A(QHSM[10]), .B(QHSM[9]), .C(CACHEPHASE), .D(n3638), .E(
        n3651), .Y(n3781) );
    zor3b U2144 ( .A(QHSM[13]), .B(QHDWNUM[0]), .C(n3781), .Y(n3782) );
    zor3b U2145 ( .A(n3652), .B(n3651), .C(n3646), .Y(n3784) );
    zao211b U2146 ( .A(n3787), .B(NXTISSTSWB), .C(n2926), .D(n3788), .Y(n3131)
         );
    zor2d U2147 ( .A(DWCNT[3]), .B(n3789), .Y(n3790) );
    zor3b U2148 ( .A(DWCNT[1]), .B(DWCNT[2]), .C(n3790), .Y(n3791) );
    zor2d U2149 ( .A(QHDWNUM[0]), .B(n3791), .Y(n3792) );
    zor3b U2150 ( .A(DWCNT[0]), .B(DWCNT[1]), .C(DWCNT[2]), .Y(n3794) );
    zor3b U2151 ( .A(n3799), .B(n3793), .C(n3790), .Y(n3801) );
    zor3b U2152 ( .A(DWCNT[1]), .B(n3799), .C(n3790), .Y(n3802) );
    zor3b U2153 ( .A(DWCNT[2]), .B(n3793), .C(n3798), .Y(n3803) );
    zor3b U2154 ( .A(n3793), .B(n3799), .C(n3798), .Y(n3804) );
    zao211b U2155 ( .A(n3354), .B(TRAN_CMD[14]), .C(n3809), .D(n3807), .Y(
        n3808) );
    zor2d U2156 ( .A(n3812), .B(n3813), .Y(n3146) );
    zor2d U2157 ( .A(n3814), .B(n3813), .Y(n3144) );
    zor3b U2158 ( .A(n3631), .B(n3104), .C(n3360), .Y(n3816) );
    zor3b U2159 ( .A(n2891), .B(n3752), .C(n3607), .Y(n3818) );
    zxo2d U2160 ( .A(n3514), .B(n3823), .Y(n3693) );
    zxo2d U2161 ( .A(n3504), .B(n3824), .Y(n3692) );
    zxo2d U2162 ( .A(n3508), .B(n3825), .Y(n3691) );
    zcx8d U2163 ( .A(n3550), .B(n3753), .C(QHSM[3]), .D(n2921), .E(n3556), .Y(
        n3830) );
    zao211b U2164 ( .A(n3787), .B(NXTISSTSWB), .C(n3833), .D(n3788), .Y(n3832)
         );
    zor3b U2165 ( .A(TRAN_CMD[6]), .B(DW2[30]), .C(n3632), .Y(n3838) );
    zoai2x4d U2166 ( .A(n3527), .B(n3512), .C(n3663), .D(n3510), .E(n3662), 
        .F(n3508), .G(n3661), .H(n3506), .Y(n3680) );
    zoai2x4d U2167 ( .A(n3660), .B(n3684), .C(n3659), .D(n3683), .E(n3658), 
        .F(n3682), .G(n3603), .H(n3681), .Y(n3845) );
    zor3b U2168 ( .A(CRCERR), .B(PIDERR), .C(RXPIDERR), .Y(n3850) );
    zan4b U2169 ( .A(n3635), .B(n3636), .C(n3634), .D(n3637), .Y(n3542) );
    zao222b U2170 ( .A(DW11[27]), .B(n3948), .C(DW10[27]), .D(n3851), .E(n3852
        ), .F(DW9[27]), .Y(n3372) );
    zao222b U2171 ( .A(DW11[26]), .B(n3745), .C(DW10[26]), .D(n3851), .E(DW9
        [26]), .F(n3852), .Y(n3374) );
    zao222b U2172 ( .A(DW11[25]), .B(n3948), .C(DW10[25]), .D(n3851), .E(DW9
        [25]), .F(n3852), .Y(n3376) );
    zao222b U2173 ( .A(DW11[24]), .B(n3745), .C(DW10[24]), .D(n3851), .E(DW9
        [24]), .F(n3852), .Y(n3378) );
    zao222b U2174 ( .A(DW11[23]), .B(n3948), .C(DW10[23]), .D(n3851), .E(DW9
        [23]), .F(n3852), .Y(n3380) );
    zao222b U2175 ( .A(DW11[22]), .B(n3745), .C(DW10[22]), .D(n3851), .E(DW9
        [22]), .F(n3852), .Y(n3382) );
    zao222b U2176 ( .A(DW11[21]), .B(n3948), .C(DW10[21]), .D(n3851), .E(DW9
        [21]), .F(n3852), .Y(n3384) );
    zao222b U2177 ( .A(DW11[20]), .B(n3745), .C(DW10[20]), .D(n3851), .E(DW9
        [20]), .F(n3852), .Y(n3386) );
    zao222b U2178 ( .A(DW11[19]), .B(n3948), .C(DW10[19]), .D(n3851), .E(DW9
        [19]), .F(n3852), .Y(n3388) );
    zao222b U2179 ( .A(DW11[18]), .B(n3745), .C(DW10[18]), .D(n3851), .E(DW9
        [18]), .F(n3852), .Y(n3390) );
    zao222b U2180 ( .A(DW11[17]), .B(n3948), .C(DW10[17]), .D(n3851), .E(DW9
        [17]), .F(n3852), .Y(n3392) );
    zao222b U2181 ( .A(DW11[16]), .B(n3745), .C(DW10[16]), .D(n3851), .E(DW9
        [16]), .F(n3852), .Y(n3394) );
    zao222b U2182 ( .A(DW11[15]), .B(n3948), .C(DW10[15]), .D(n3851), .E(DW9
        [15]), .F(n3852), .Y(n3396) );
    zao222b U2183 ( .A(DW11[14]), .B(n3745), .C(DW10[14]), .D(n3851), .E(DW9
        [14]), .F(n3852), .Y(n3398) );
    zao222b U2184 ( .A(DW11[13]), .B(n3948), .C(DW10[13]), .D(n3851), .E(DW9
        [13]), .F(n3852), .Y(n3400) );
    zao222b U2185 ( .A(DW11[12]), .B(n3745), .C(DW10[12]), .D(n3851), .E(DW9
        [12]), .F(n3852), .Y(n3402) );
    zao222b U2186 ( .A(DW11[31]), .B(n3948), .C(DW10[31]), .D(n3851), .E(DW9
        [31]), .F(n3852), .Y(n3364) );
    zao222b U2187 ( .A(DW11[30]), .B(n3745), .C(DW10[30]), .D(n3851), .E(DW9
        [30]), .F(n3852), .Y(n3366) );
    zao222b U2188 ( .A(DW11[29]), .B(n3948), .C(DW10[29]), .D(n3851), .E(DW9
        [29]), .F(n3852), .Y(n3368) );
    zao222b U2189 ( .A(DW11[28]), .B(n3948), .C(DW10[28]), .D(n3851), .E(DW9
        [28]), .F(n3852), .Y(n3370) );
    zor3b U2190 ( .A(n3552), .B(n3555), .C(QTDHALT), .Y(n3833) );
    zcx8d U2191 ( .A(EHCI_MAC_EOT), .B(n3778), .C(n3490), .D(IMMEDRETRY), .E(
        n3566), .Y(n3779) );
    zor4b U2192 ( .A(DW6[7]), .B(DW6[6]), .C(n3577), .D(n3650), .Y(n3570) );
    zao222b U2193 ( .A(QHSM[9]), .B(QHSM[11]), .C(QHSM[13]), .D(n2930), .E(
        n3573), .F(QHCIMWR), .Y(n3853) );
    zor3b U2194 ( .A(n3835), .B(n3859), .C(n3860), .Y(n3088) );
    zao211b U2195 ( .A(PCIEND), .B(n3861), .C(GEN_PERR), .D(n3585), .Y(n3860)
         );
    zao222b U2196 ( .A(QHSM[4]), .B(QHSM[1]), .C(QHSM[0]), .D(n3586), .E(n3651
        ), .F(n3646), .Y(n3859) );
    zao222b U2197 ( .A(n3863), .B(DW11[9]), .C(DW7[9]), .D(n3944), .E(DW3[9]), 
        .F(n3946), .Y(n3272) );
    zao222b U2198 ( .A(DW11[8]), .B(n3942), .C(DW7[8]), .D(n3864), .E(DW3[8]), 
        .F(n3865), .Y(n3270) );
    zao222b U2199 ( .A(DW11[7]), .B(n3863), .C(DW7[7]), .D(n3944), .E(DW3[7]), 
        .F(n3946), .Y(n3268) );
    zao222b U2200 ( .A(DW11[6]), .B(n3942), .C(DW7[6]), .D(n3943), .E(DW3[6]), 
        .F(n3945), .Y(n3266) );
    zao222b U2201 ( .A(DW11[5]), .B(n3863), .C(DW7[5]), .D(n3864), .E(DW3[5]), 
        .F(n3865), .Y(n3264) );
    zao211b U2202 ( .A(DW4[4]), .B(n3947), .C(n3875), .D(n3876), .Y(n3261) );
    zao222b U2203 ( .A(DW11[4]), .B(n3942), .C(DW7[4]), .D(n3943), .E(DW3[4]), 
        .F(n3945), .Y(n3262) );
    zao222b U2204 ( .A(n3942), .B(DW11[31]), .C(DW7[31]), .D(n3944), .E(DW3
        [31]), .F(n3946), .Y(n3316) );
    zao222b U2205 ( .A(n3863), .B(DW11[30]), .C(DW7[30]), .D(n3864), .E(DW3
        [30]), .F(n3865), .Y(n3314) );
    zao211b U2206 ( .A(DW4[3]), .B(n3874), .C(n3879), .D(n3880), .Y(n3259) );
    zao222b U2207 ( .A(DW11[3]), .B(n3863), .C(DW7[3]), .D(n3943), .E(DW3[3]), 
        .F(n3945), .Y(n3260) );
    zao222b U2208 ( .A(n3942), .B(DW11[29]), .C(DW7[29]), .D(n3944), .E(DW3
        [29]), .F(n3946), .Y(n3312) );
    zao222b U2209 ( .A(n3863), .B(DW11[28]), .C(DW7[28]), .D(n3864), .E(DW3
        [28]), .F(n3865), .Y(n3310) );
    zao222b U2210 ( .A(n3942), .B(DW11[27]), .C(DW7[27]), .D(n3943), .E(DW3
        [27]), .F(n3945), .Y(n3308) );
    zao222b U2211 ( .A(n3863), .B(DW11[26]), .C(DW7[26]), .D(n3944), .E(DW3
        [26]), .F(n3946), .Y(n3306) );
    zao222b U2212 ( .A(n3942), .B(DW11[25]), .C(DW7[25]), .D(n3864), .E(DW3
        [25]), .F(n3865), .Y(n3304) );
    zao222b U2213 ( .A(n3863), .B(DW11[24]), .C(DW7[24]), .D(n3943), .E(DW3
        [24]), .F(n3945), .Y(n3302) );
    zao222b U2214 ( .A(n3942), .B(DW11[23]), .C(DW7[23]), .D(n3944), .E(DW3
        [23]), .F(n3946), .Y(n3300) );
    zao222b U2215 ( .A(n3863), .B(DW11[22]), .C(DW7[22]), .D(n3864), .E(DW3
        [22]), .F(n3865), .Y(n3298) );
    zao222b U2216 ( .A(n3942), .B(DW11[21]), .C(DW7[21]), .D(n3943), .E(DW3
        [21]), .F(n3945), .Y(n3296) );
    zao222b U2217 ( .A(n3863), .B(DW11[20]), .C(DW7[20]), .D(n3944), .E(DW3
        [20]), .F(n3946), .Y(n3294) );
    zao211b U2218 ( .A(DW4[2]), .B(n3947), .C(n3891), .D(n3892), .Y(n3257) );
    zao222b U2219 ( .A(DW11[2]), .B(n3942), .C(DW7[2]), .D(n3864), .E(DW3[2]), 
        .F(n3865), .Y(n3258) );
    zao222b U2220 ( .A(n3942), .B(DW11[19]), .C(DW7[19]), .D(n3943), .E(DW3
        [19]), .F(n3945), .Y(n3292) );
    zao222b U2221 ( .A(n3863), .B(DW11[18]), .C(DW7[18]), .D(n3944), .E(DW3
        [18]), .F(n3946), .Y(n3290) );
    zao222b U2222 ( .A(n3942), .B(DW11[17]), .C(DW7[17]), .D(n3864), .E(DW3
        [17]), .F(n3865), .Y(n3288) );
    zao222b U2223 ( .A(n3863), .B(DW11[16]), .C(DW7[16]), .D(n3944), .E(DW3
        [16]), .F(n3945), .Y(n3286) );
    zao222b U2224 ( .A(n3942), .B(DW11[15]), .C(DW7[15]), .D(n3943), .E(DW3
        [15]), .F(n3946), .Y(n3284) );
    zao222b U2225 ( .A(n3863), .B(DW11[14]), .C(DW7[14]), .D(n3864), .E(DW3
        [14]), .F(n3865), .Y(n3282) );
    zoai2x4d U2226 ( .A(n3803), .B(n3214), .C(n3415), .D(n3951), .E(n3416), 
        .F(n3953), .G(n3417), .H(n3955), .Y(n3898) );
    zao222b U2227 ( .A(n3942), .B(DW11[13]), .C(DW7[13]), .D(n3943), .E(DW3
        [13]), .F(n3945), .Y(n3280) );
    zao222b U2228 ( .A(n3863), .B(DW11[12]), .C(DW7[12]), .D(n3944), .E(DW3
        [12]), .F(n3946), .Y(n3278) );
    zao222b U2229 ( .A(DW11[11]), .B(n3863), .C(DW7[11]), .D(n3864), .E(DW3
        [11]), .F(n3865), .Y(n3276) );
    zao222b U2230 ( .A(DW11[10]), .B(n3942), .C(DW7[10]), .D(n3943), .E(DW3
        [10]), .F(n3945), .Y(n3274) );
    zao211b U2231 ( .A(DW4[1]), .B(n3874), .C(n3903), .D(n3904), .Y(n3255) );
    zao222b U2232 ( .A(DW11[1]), .B(n3863), .C(DW7[1]), .D(n3944), .E(DW3[1]), 
        .F(n3946), .Y(n3256) );
    zao222b U2233 ( .A(DW11[0]), .B(n3942), .C(DW7[0]), .D(n3864), .E(DW3[0]), 
        .F(n3865), .Y(n3254) );
    zor6b U2234 ( .A(MAXLEN[7]), .B(MAXLEN[6]), .C(MAXLEN[5]), .D(MAXLEN[10]), 
        .E(MAXLEN[9]), .F(MAXLEN[8]), .Y(n3593) );
    zor3b U2235 ( .A(n2926), .B(n3776), .C(n3091), .Y(n3109) );
    zor3b U2236 ( .A(DW6[9]), .B(n3699), .C(n3748), .Y(n3547) );
    zor4b U2237 ( .A(n3610), .B(n2893), .C(n3129), .D(n3753), .Y(n3613) );
    zor4b U2238 ( .A(n3559), .B(n3523), .C(n2868), .D(n3520), .Y(n3564) );
    zivh U2239 ( .A(n3633), .Y(n3358) );
    zor2d U2240 ( .A(n3349), .B(UP_DW8[2]), .Y(n3825) );
    zor2d U2241 ( .A(n3351), .B(UP_DW8[4]), .Y(n3824) );
    zor2d U2242 ( .A(n3354), .B(UP_DW8[7]), .Y(n3823) );
    zor2d U2243 ( .A(n3352), .B(UP_DW8[5]), .Y(n3822) );
    zor2d U2244 ( .A(n3353), .B(UP_DW8[6]), .Y(n3821) );
    zor2d U2245 ( .A(n3350), .B(UP_DW8[3]), .Y(n3820) );
    zor2d U2246 ( .A(n3348), .B(UP_DW8[1]), .Y(n3819) );
    zao211b U2247 ( .A(TMOUT), .B(n3920), .C(n3850), .D(n3529), .Y(n3533) );
    zao211b U2248 ( .A(RXPIDERR), .B(n3358), .C(n3774), .D(n3753), .Y(n3536)
         );
    zor3b U2249 ( .A(n2892), .B(n3627), .C(n2921), .Y(n3545) );
    zor3b U2250 ( .A(n3566), .B(n3491), .C(n3553), .Y(n3551) );
    zor4b U2251 ( .A(n3518), .B(n3678), .C(n2868), .D(n3517), .Y(n3558) );
    zor3b U2252 ( .A(n3642), .B(n3523), .C(n3557), .Y(n3780) );
    zor2d U2253 ( .A(n3642), .B(n2889), .Y(n3581) );
    zor3b U2254 ( .A(n3626), .B(n3518), .C(n3517), .Y(n3560) );
    zor4b U2255 ( .A(n3572), .B(n3853), .C(n3854), .D(n3584), .Y(n3924) );
    zao211b U2256 ( .A(n3909), .B(n3578), .C(n2876), .D(n3574), .Y(n3861) );
    zor4b U2257 ( .A(DW6[6]), .B(n3133), .C(n2888), .D(n3576), .Y(n3087) );
    zao32d U2258 ( .A(n2925), .B(n3793), .C(n3919), .D(n3908), .E(QHDWNUM[0]), 
        .Y(n3864) );
    zao22d U2259 ( .A(QHDWNUM[3]), .B(n3907), .C(DWCNT[3]), .D(n3794), .Y(
        n3865) );
    zao32d U2260 ( .A(n2924), .B(n3799), .C(n3918), .D(n3907), .E(n3797), .Y(
        n3252) );
    zor3b U2261 ( .A(QHSM[7]), .B(QHSM[8]), .C(n3594), .Y(n3101) );
    zoai21d U2262 ( .A(n3922), .B(n3360), .C(n3766), .Y(n3331) );
    zao222b U2263 ( .A(OVERWBOFFSET_P2070_9), .B(TRAN_CMD[9]), .C(n3609), .D(
        TRAN_CMD[81]), .E(OVERWBOFFSET_P2090_9), .F(n3608), .Y(n3342) );
    zao222b U2264 ( .A(OVERWBOFFSET_P2070_8), .B(TRAN_CMD[9]), .C(TRAN_CMD[80]
        ), .D(n3609), .E(OVERWBOFFSET_P2090_8), .F(n3608), .Y(n3341) );
    zao222b U2265 ( .A(OVERWBOFFSET_P2070_7), .B(UP_DW6[8]), .C(TRAN_CMD[79]), 
        .D(n3609), .E(OVERWBOFFSET_P2090_7), .F(n3608), .Y(n3340) );
    zao222b U2266 ( .A(OVERWBOFFSET_P2070_6), .B(TRAN_CMD[9]), .C(TRAN_CMD[78]
        ), .D(n3609), .E(OVERWBOFFSET_P2090_6), .F(n3608), .Y(n3339) );
    zao222b U2267 ( .A(OVERWBOFFSET_P2070_5), .B(UP_DW6[8]), .C(TRAN_CMD[77]), 
        .D(n3609), .E(OVERWBOFFSET_P2090_5), .F(n3608), .Y(n3338) );
    zao222b U2268 ( .A(OVERWBOFFSET_P2070_4), .B(TRAN_CMD[9]), .C(TRAN_CMD[76]
        ), .D(n3609), .E(OVERWBOFFSET_P2090_4), .F(n3608), .Y(n3337) );
    zao222b U2269 ( .A(OVERWBOFFSET_P2070_3), .B(TRAN_CMD[9]), .C(TRAN_CMD[75]
        ), .D(n3609), .E(OVERWBOFFSET_P2090_3), .F(n3608), .Y(n3336) );
    zao222b U2270 ( .A(OVERWBOFFSET_P2070_2), .B(TRAN_CMD[9]), .C(TRAN_CMD[74]
        ), .D(n3609), .E(OVERWBOFFSET_P2090_2), .F(n3608), .Y(n3335) );
    zao222b U2271 ( .A(OVERWBOFFSET_P2070_11), .B(TRAN_CMD[9]), .C(TRAN_CMD
        [83]), .D(n3609), .E(OVERWBOFFSET_P2090_11), .F(n3608), .Y(n3344) );
    zao222b U2272 ( .A(OVERWBOFFSET_P2070_10), .B(TRAN_CMD[9]), .C(TRAN_CMD
        [82]), .D(n3609), .E(OVERWBOFFSET_P2090_10), .F(n3608), .Y(n3343) );
    zao222b U2273 ( .A(OVERWBOFFSET_P2070_1), .B(TRAN_CMD[9]), .C(TRAN_CMD[73]
        ), .D(n3609), .E(OVERWBOFFSET_P2090_1), .F(n3608), .Y(n3334) );
    zao222b U2274 ( .A(OVERWBOFFSET_P2070_0), .B(UP_DW6[8]), .C(TRAN_CMD[72]), 
        .D(n3609), .E(OVERWBOFFSET_P2090_0), .F(n3608), .Y(n3333) );
    zor2d U2275 ( .A(n3345), .B(n2872), .Y(n3347) );
    zor3b U2276 ( .A(QHSM[2]), .B(CACHE_MODIFY), .C(PHASENXT_resultwb), .Y(
        n3317) );
    zor3b U2277 ( .A(TRAN_CMD[14]), .B(n3764), .C(QHDWNUM[2]), .Y(n3616) );
    zmux21ld U2278 ( .A(n3126), .B(n3530), .S(n2932), .Y(n3319) );
    zor4b U2279 ( .A(n3590), .B(n2881), .C(n2908), .D(n3619), .Y(n3844) );
    zor2d U2280 ( .A(n3814), .B(n3813), .Y(n3929) );
    zor2d U2281 ( .A(n3814), .B(n3813), .Y(n3930) );
    zor2d U2282 ( .A(n3812), .B(n3813), .Y(n3931) );
    zor2d U2283 ( .A(n3812), .B(n3813), .Y(n3932) );
    zao32d U2284 ( .A(DWCNT[1]), .B(n3799), .C(n3918), .D(n3907), .E(n3797), 
        .Y(n3933) );
    zao32d U2285 ( .A(n2924), .B(n3799), .C(n3918), .D(n3907), .E(n3797), .Y(
        n3934) );
    zor3b U2286 ( .A(n3746), .B(n3747), .C(n3745), .Y(n3935) );
    zor3b U2287 ( .A(n3746), .B(n3747), .C(n3948), .Y(n3936) );
    zor3b U2288 ( .A(n3747), .B(n3745), .C(n3630), .Y(n3937) );
    zor3b U2289 ( .A(n3747), .B(n3948), .C(n3630), .Y(n3938) );
    zor3b U2290 ( .A(n3746), .B(n3745), .C(n3628), .Y(n3939) );
    zor3b U2291 ( .A(n3746), .B(n3948), .C(n3628), .Y(n3940) );
    zao32d U2292 ( .A(DWCNT[2]), .B(n3793), .C(n3919), .D(n3908), .E(QHDWNUM
        [0]), .Y(n3943) );
    zao32d U2293 ( .A(n2925), .B(n3793), .C(n3919), .D(n3908), .E(QHDWNUM[0]), 
        .Y(n3944) );
    zao22d U2294 ( .A(QHDWNUM[3]), .B(n3907), .C(DWCNT[3]), .D(n3794), .Y(
        n3945) );
    zao22d U2295 ( .A(QHDWNUM[3]), .B(n3907), .C(DWCNT[3]), .D(n3794), .Y(
        n3946) );
    zor3b U2296 ( .A(DWCNT[2]), .B(n3793), .C(n3798), .Y(n3949) );
    zor3b U2297 ( .A(DWCNT[2]), .B(n3793), .C(n3798), .Y(n3950) );
    zor3b U2298 ( .A(DWCNT[1]), .B(n3799), .C(n3790), .Y(n3951) );
    zor3b U2299 ( .A(DWCNT[1]), .B(n3799), .C(n3790), .Y(n3952) );
    zor3b U2300 ( .A(n3793), .B(n3799), .C(n3798), .Y(n3953) );
    zor3b U2301 ( .A(n3793), .B(n3799), .C(n3798), .Y(n3954) );
    zor3b U2302 ( .A(n3799), .B(n3793), .C(n3790), .Y(n3955) );
    zor3b U2303 ( .A(n3799), .B(n3793), .C(n3790), .Y(n3956) );
endmodule


module PERIODIC_MUX ( TD_CACHE_EN1, TD_CACHE_EN2, EXEITD1, EXEITD2, EXEQH1, 
    EXEQH2, EXESITD1, EXESITD2, DWNUM, IDWNUM1, QHDWNUM1, SIDWNUM1, IDWNUM2, 
    QHDWNUM2, SIDWNUM2, IDWOFFSET1, QHDWOFFSET1, SIDWOFFSET1, IDWOFFSET2, 
    QHDWOFFSET2, SIDWOFFSET2, EDWNUM, DWOFFSET, EDWOFFSET, QUP_DW1_3, 
    SIUP_DW1_3, UP_DW1_3, QUP_DW2_3, SIUP_DW2_3, UP_DW2_3, QUP_LDW1_3, 
    SIUP_LDW1_3, UP_LDW1_3, QUP_LDW2_3, SIUP_LDW2_3, UP_LDW2_3, QCACHEPHASE1, 
    QCACHEPHASE2, SICACHEPHASE1, SICACHEPHASE2, CACHEPHASE1, CACHEPHASE2, 
    EHCI_MAC_EOT, IHCIREQ1, IHCIREQ2, QHCIREQ1, QHCIREQ2, SIHCIREQ1, SIHCIREQ2, 
    TDHCIREQ1, TDHCIREQ2, TDHCIGNT1, TDHCIGNT2, IMWR1, QHMWR1, SIMWR1, IMWR2, 
    QHMWR2, SIMWR2, HCIMWR, PCIEND, IPCIEND1, IPCIEND2, QPCIEND1, QPCIEND2, 
    SIPCIEND1, SIPCIEND2, TD_ACT1, TD_ACT2, ITD_ACT1, ITD_ACT2, QH_ACT1, 
    QH_ACT2, SITD_ACT1, SITD_ACT2, ITD_MAC_EOT1, ITD_MAC_EOT2, QH_MAC_EOT1, 
    QH_MAC_EOT2, SITD_MAC_EOT1, SITD_MAC_EOT2, PARSEITDEND1, PARSEITDEND2, 
    PARSEQHEND1, PARSEQHEND2, PARSESITDEND1, PARSESITDEND2, PARSETDEND1, 
    PARSETDEND2, ITDPARSING1, ITDPARSING2, QHPARSING1, QHPARSING2, 
    SITDPARSING1, SITDPARSING2, TDPARSING1, TDPARSING2, TD_PARSE_GO1, 
    TD_PARSE_GO2, ITD_PARSE_GO1, ITD_PARSE_GO2, QH_PARSE_GO1, QH_PARSE_GO2, 
    SITD_PARSE_GO1, SITD_PARSE_GO2, ICACHE_INVALID1, ICACHE_INVALID2, 
    QCACHE_INVALID1, QCACHE_INVALID2, SICACHE_INVALID1, SICACHE_INVALID2, 
    CACHE_INVALID1, CACHE_INVALID2, ICMDSTART_REQ1, ICMDSTART_REQ2, 
    QCMDSTART_REQ1, QCMDSTART_REQ2, SICMDSTART_REQ1, SICMDSTART_REQ2, 
    PER_CMDSTART_REQ1, PER_CMDSTART_REQ2, PER_CMDSTART1, PER_CMDSTART2, 
    ICMDSTART1, ICMDSTART2, QCMDSTART1, QCMDSTART2, SICMDSTART1, SICMDSTART2, 
    ITRAN_CMD1, ITRAN_CMD2, QTRAN_CMD1, QTRAN_CMD2, SITRAN_CMD1, SITRAN_CMD2, 
    TRAN_CMD1, TRAN_CMD2, IBUI_GO1, IBUI_GO2, QBUI_GO1, QBUI_GO2, SIBUI_GO1, 
    SIBUI_GO2, BUI_GO1, BUI_GO2, IRXERR1, IRXERR2, QRXERR1, QRXERR2, SIRXERR1, 
    SIRXERR2, RXERR1, RXERR2, IEOT1, IEOT2, QEOT1, QEOT2, SIEOT1, SIEOT2, EOT1, 
    EOT2, USBDMA_SEL, CRCERR, BABBLE, PIDERR, TMOUT, TOGMATCH, RXNAK, RXNYET, 
    RXSTALL, RXACK, RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXPIDERR, SPD, ACTLEN, 
    CRCERR1, BABBLE1, PIDERR1, TMOUT1, TOGMATCH1, RXNAK1, RXNYET1, RXSTALL1, 
    RXACK1, RXDATA01, RXDATA11, RXDATA21, RXMDATA1, RXPIDERR1, SPD1, ACTLEN1, 
    CRCERR2, BABBLE2, PIDERR2, TMOUT2, TOGMATCH2, RXNAK2, RXNYET2, RXSTALL2, 
    RXACK2, RXDATA02, RXDATA12, RXDATA22, RXMDATA2, RXPIDERR2, SPD2, ACTLEN2
     );
input  [3:0] DWNUM;
input  [3:0] IDWNUM1;
input  [3:0] SIDWNUM1;
input  [31:0] QUP_DW1_3;
input  [104:0] QTRAN_CMD2;
input  [3:0] IDWOFFSET1;
input  [104:0] SITRAN_CMD1;
output [104:0] TRAN_CMD2;
input  [3:0] QHDWNUM1;
input  [3:0] SIDWOFFSET2;
input  [3:0] DWOFFSET;
input  [104:0] ITRAN_CMD2;
output [10:0] ACTLEN1;
output [31:0] UP_DW1_3;
input  [4:0] USBDMA_SEL;
input  [3:0] IDWNUM2;
input  [3:0] SIDWNUM2;
input  [3:0] QHDWOFFSET2;
output [3:0] EDWNUM;
input  [31:0] SIUP_DW1_3;
input  [104:0] QTRAN_CMD1;
input  [3:0] IDWOFFSET2;
output [3:0] EDWOFFSET;
input  [31:0] SIUP_DW2_3;
output [31:0] UP_DW2_3;
input  [104:0] SITRAN_CMD2;
output [104:0] TRAN_CMD1;
input  [10:0] ACTLEN;
input  [3:0] QHDWNUM2;
input  [3:0] SIDWOFFSET1;
input  [31:0] QUP_DW2_3;
input  [104:0] ITRAN_CMD1;
output [10:0] ACTLEN2;
input  [3:0] QHDWOFFSET1;
input  TD_CACHE_EN1, TD_CACHE_EN2, EXEITD1, EXEITD2, EXEQH1, EXEQH2, EXESITD1, 
    EXESITD2, QUP_LDW1_3, SIUP_LDW1_3, QUP_LDW2_3, SIUP_LDW2_3, QCACHEPHASE1, 
    QCACHEPHASE2, SICACHEPHASE1, SICACHEPHASE2, EHCI_MAC_EOT, IHCIREQ1, 
    IHCIREQ2, QHCIREQ1, QHCIREQ2, SIHCIREQ1, SIHCIREQ2, TDHCIGNT1, TDHCIGNT2, 
    IMWR1, QHMWR1, SIMWR1, IMWR2, QHMWR2, SIMWR2, PCIEND, TD_ACT1, TD_ACT2, 
    PARSEITDEND1, PARSEITDEND2, PARSEQHEND1, PARSEQHEND2, PARSESITDEND1, 
    PARSESITDEND2, ITDPARSING1, ITDPARSING2, QHPARSING1, QHPARSING2, 
    SITDPARSING1, SITDPARSING2, TD_PARSE_GO1, TD_PARSE_GO2, ICACHE_INVALID1, 
    ICACHE_INVALID2, QCACHE_INVALID1, QCACHE_INVALID2, SICACHE_INVALID1, 
    SICACHE_INVALID2, ICMDSTART_REQ1, ICMDSTART_REQ2, QCMDSTART_REQ1, 
    QCMDSTART_REQ2, SICMDSTART_REQ1, SICMDSTART_REQ2, PER_CMDSTART1, 
    PER_CMDSTART2, IBUI_GO1, IBUI_GO2, QBUI_GO1, QBUI_GO2, SIBUI_GO1, 
    SIBUI_GO2, IRXERR1, IRXERR2, QRXERR1, QRXERR2, SIRXERR1, SIRXERR2, IEOT1, 
    IEOT2, QEOT1, QEOT2, SIEOT1, SIEOT2, CRCERR, BABBLE, PIDERR, TMOUT, 
    TOGMATCH, RXNAK, RXNYET, RXSTALL, RXACK, RXDATA0, RXDATA1, RXDATA2, 
    RXMDATA, RXPIDERR, SPD;
output UP_LDW1_3, UP_LDW2_3, CACHEPHASE1, CACHEPHASE2, TDHCIREQ1, TDHCIREQ2, 
    HCIMWR, IPCIEND1, IPCIEND2, QPCIEND1, QPCIEND2, SIPCIEND1, SIPCIEND2, 
    ITD_ACT1, ITD_ACT2, QH_ACT1, QH_ACT2, SITD_ACT1, SITD_ACT2, ITD_MAC_EOT1, 
    ITD_MAC_EOT2, QH_MAC_EOT1, QH_MAC_EOT2, SITD_MAC_EOT1, SITD_MAC_EOT2, 
    PARSETDEND1, PARSETDEND2, TDPARSING1, TDPARSING2, ITD_PARSE_GO1, 
    ITD_PARSE_GO2, QH_PARSE_GO1, QH_PARSE_GO2, SITD_PARSE_GO1, SITD_PARSE_GO2, 
    CACHE_INVALID1, CACHE_INVALID2, PER_CMDSTART_REQ1, PER_CMDSTART_REQ2, 
    ICMDSTART1, ICMDSTART2, QCMDSTART1, QCMDSTART2, SICMDSTART1, SICMDSTART2, 
    BUI_GO1, BUI_GO2, RXERR1, RXERR2, EOT1, EOT2, CRCERR1, BABBLE1, PIDERR1, 
    TMOUT1, TOGMATCH1, RXNAK1, RXNYET1, RXSTALL1, RXACK1, RXDATA01, RXDATA11, 
    RXDATA21, RXMDATA1, RXPIDERR1, SPD1, CRCERR2, BABBLE2, PIDERR2, TMOUT2, 
    TOGMATCH2, RXNAK2, RXNYET2, RXSTALL2, RXACK2, RXDATA02, RXDATA12, RXDATA22, 
    RXMDATA2, RXPIDERR2, SPD2;
    wire n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
        n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
        n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
        n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
        n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
        n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
        n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
        n1679, n1680, n1681, n1682;
    zivd U67 ( .A(n1613), .Y(n1640) );
    zivd U68 ( .A(n1652), .Y(n1655) );
    zivd U69 ( .A(n1647), .Y(n1650) );
    zivd U70 ( .A(n1652), .Y(n1653) );
    zivd U71 ( .A(n1647), .Y(n1648) );
    zivd U72 ( .A(n1609), .Y(n1644) );
    zivd U73 ( .A(n1611), .Y(n1641) );
    zivd U74 ( .A(n1615), .Y(n1635) );
    ziv11d U75 ( .A(n1678), .Y(n1609), .Z(n1610) );
    zinr2b U76 ( .A(EXESITD2), .B(n1639), .Y(n1678) );
    ziv11d U77 ( .A(n1677), .Y(n1611), .Z(n1612) );
    zinr2b U78 ( .A(EXESITD1), .B(n1637), .Y(n1677) );
    ziv11d U79 ( .A(EXEITD2), .Y(n1613), .Z(n1614) );
    ziv11d U80 ( .A(EXEITD1), .Y(n1615), .Z(n1616) );
    zivd U81 ( .A(n1647), .Y(n1618) );
    zivd U82 ( .A(n1647), .Y(n1617) );
    zivd U83 ( .A(n1647), .Y(n1651) );
    zivd U84 ( .A(n1647), .Y(n1649) );
    zivd U85 ( .A(n1609), .Y(n1620) );
    zivd U86 ( .A(n1609), .Y(n1619) );
    zivd U87 ( .A(n1609), .Y(n1646) );
    zivd U88 ( .A(n1609), .Y(n1645) );
    zivd U89 ( .A(n1652), .Y(n1622) );
    zivd U90 ( .A(n1652), .Y(n1621) );
    zivd U91 ( .A(n1652), .Y(n1656) );
    zivd U92 ( .A(n1652), .Y(n1654) );
    zivd U93 ( .A(n1611), .Y(n1624) );
    zivd U94 ( .A(n1611), .Y(n1623) );
    zivd U95 ( .A(n1611), .Y(n1643) );
    zivd U96 ( .A(n1611), .Y(n1642) );
    zivd U97 ( .A(n1613), .Y(n1626) );
    zivd U98 ( .A(n1613), .Y(n1625) );
    zivd U99 ( .A(n1613), .Y(n1639) );
    zivd U100 ( .A(n1613), .Y(n1638) );
    zivd U101 ( .A(n1615), .Y(n1628) );
    zivd U102 ( .A(n1615), .Y(n1627) );
    zivd U103 ( .A(n1615), .Y(n1636) );
    zivd U104 ( .A(n1615), .Y(n1637) );
    zbfd U105 ( .A(USBDMA_SEL[1]), .Y(n1629) );
    zbfd U106 ( .A(USBDMA_SEL[0]), .Y(n1630) );
    zbfd U107 ( .A(EXEQH2), .Y(n1631) );
    zbfd U108 ( .A(EXEQH2), .Y(n1632) );
    zbfd U109 ( .A(EXEQH1), .Y(n1633) );
    zbfd U110 ( .A(EXEQH1), .Y(n1634) );
    zor2b U111 ( .A(n1635), .B(EXESITD1), .Y(n1647) );
    zor2b U112 ( .A(n1625), .B(EXESITD2), .Y(n1652) );
    zao222b U113 ( .A(n1657), .B(n1658), .C(DWNUM[0]), .D(n1659), .E(TDHCIGNT1
        ), .F(n1660), .Y(EDWNUM[0]) );
    zao222b U114 ( .A(n1657), .B(n1661), .C(DWNUM[1]), .D(n1659), .E(TDHCIGNT1
        ), .F(n1662), .Y(EDWNUM[1]) );
    zao222b U115 ( .A(n1657), .B(n1663), .C(DWNUM[2]), .D(n1659), .E(TDHCIGNT1
        ), .F(n1664), .Y(EDWNUM[2]) );
    zao222b U116 ( .A(n1657), .B(n1665), .C(DWNUM[3]), .D(n1659), .E(TDHCIGNT1
        ), .F(n1666), .Y(EDWNUM[3]) );
    zan2b U117 ( .A(CRCERR), .B(n1630), .Y(CRCERR1) );
    zan2b U118 ( .A(BABBLE), .B(n1630), .Y(BABBLE1) );
    zan2b U119 ( .A(PIDERR), .B(n1630), .Y(PIDERR1) );
    zan2b U120 ( .A(TMOUT), .B(n1630), .Y(TMOUT1) );
    zan2b U121 ( .A(n1630), .B(TOGMATCH), .Y(TOGMATCH1) );
    zan2b U122 ( .A(RXNAK), .B(n1630), .Y(RXNAK1) );
    zan2b U123 ( .A(RXNYET), .B(USBDMA_SEL[0]), .Y(RXNYET1) );
    zan2b U124 ( .A(RXSTALL), .B(USBDMA_SEL[0]), .Y(RXSTALL1) );
    zan2b U125 ( .A(RXACK), .B(USBDMA_SEL[0]), .Y(RXACK1) );
    zan2b U126 ( .A(RXDATA0), .B(USBDMA_SEL[0]), .Y(RXDATA01) );
    zan2b U127 ( .A(RXDATA1), .B(n1630), .Y(RXDATA11) );
    zan2b U128 ( .A(RXDATA2), .B(n1630), .Y(RXDATA21) );
    zan2b U129 ( .A(RXMDATA), .B(USBDMA_SEL[0]), .Y(RXMDATA1) );
    zan2b U130 ( .A(RXPIDERR), .B(n1630), .Y(RXPIDERR1) );
    zan2b U131 ( .A(SPD), .B(n1630), .Y(SPD1) );
    zan2b U132 ( .A(ACTLEN[10]), .B(USBDMA_SEL[0]), .Y(ACTLEN1[10]) );
    zan2b U133 ( .A(ACTLEN[9]), .B(n1630), .Y(ACTLEN1[9]) );
    zan2b U134 ( .A(ACTLEN[8]), .B(USBDMA_SEL[0]), .Y(ACTLEN1[8]) );
    zan2b U135 ( .A(ACTLEN[7]), .B(USBDMA_SEL[0]), .Y(ACTLEN1[7]) );
    zan2b U136 ( .A(ACTLEN[6]), .B(n1630), .Y(ACTLEN1[6]) );
    zan2b U137 ( .A(ACTLEN[5]), .B(n1630), .Y(ACTLEN1[5]) );
    zan2b U138 ( .A(ACTLEN[4]), .B(n1630), .Y(ACTLEN1[4]) );
    zan2b U139 ( .A(ACTLEN[3]), .B(n1630), .Y(ACTLEN1[3]) );
    zan2b U140 ( .A(ACTLEN[2]), .B(n1630), .Y(ACTLEN1[2]) );
    zan2b U141 ( .A(ACTLEN[1]), .B(n1630), .Y(ACTLEN1[1]) );
    zan2b U142 ( .A(ACTLEN[0]), .B(n1630), .Y(ACTLEN1[0]) );
    zao222b U143 ( .A(n1667), .B(n1668), .C(DWOFFSET[0]), .D(n1669), .E(
        TD_CACHE_EN1), .F(n1670), .Y(EDWOFFSET[0]) );
    zao222b U144 ( .A(n1667), .B(n1671), .C(DWOFFSET[1]), .D(n1669), .E(
        TD_CACHE_EN1), .F(n1672), .Y(EDWOFFSET[1]) );
    zao222b U145 ( .A(n1667), .B(n1673), .C(DWOFFSET[2]), .D(n1669), .E(
        TD_CACHE_EN1), .F(n1674), .Y(EDWOFFSET[2]) );
    zao222b U146 ( .A(n1667), .B(n1675), .C(DWOFFSET[3]), .D(n1669), .E(
        TD_CACHE_EN1), .F(n1676), .Y(EDWOFFSET[3]) );
    zao222b U147 ( .A(SITRAN_CMD1[0]), .B(n1624), .C(QTRAN_CMD1[0]), .D(n1649), 
        .E(ITRAN_CMD1[0]), .F(n1636), .Y(TRAN_CMD1[0]) );
    zao222b U148 ( .A(SITRAN_CMD1[1]), .B(n1624), .C(QTRAN_CMD1[1]), .D(n1651), 
        .E(ITRAN_CMD1[1]), .F(n1635), .Y(TRAN_CMD1[1]) );
    zao222b U149 ( .A(SITRAN_CMD1[2]), .B(n1641), .C(QTRAN_CMD1[2]), .D(n1650), 
        .E(ITRAN_CMD1[2]), .F(n1616), .Y(TRAN_CMD1[2]) );
    zao222b U150 ( .A(SITRAN_CMD1[3]), .B(n1623), .C(QTRAN_CMD1[3]), .D(n1618), 
        .E(ITRAN_CMD1[3]), .F(n1628), .Y(TRAN_CMD1[3]) );
    zao222b U151 ( .A(SITRAN_CMD1[4]), .B(n1643), .C(QTRAN_CMD1[4]), .D(n1649), 
        .E(ITRAN_CMD1[4]), .F(n1636), .Y(TRAN_CMD1[4]) );
    zao222b U152 ( .A(SITRAN_CMD1[5]), .B(n1623), .C(QTRAN_CMD1[5]), .D(n1618), 
        .E(ITRAN_CMD1[5]), .F(n1628), .Y(TRAN_CMD1[5]) );
    zao222b U153 ( .A(SITRAN_CMD1[6]), .B(n1612), .C(QTRAN_CMD1[6]), .D(n1651), 
        .E(ITRAN_CMD1[6]), .F(n1635), .Y(TRAN_CMD1[6]) );
    zao222b U154 ( .A(SITRAN_CMD1[7]), .B(n1642), .C(QTRAN_CMD1[7]), .D(n1648), 
        .E(ITRAN_CMD1[7]), .F(n1616), .Y(TRAN_CMD1[7]) );
    zao222b U155 ( .A(SITRAN_CMD1[8]), .B(n1641), .C(QTRAN_CMD1[8]), .D(n1651), 
        .E(ITRAN_CMD1[8]), .F(n1635), .Y(TRAN_CMD1[8]) );
    zao222b U156 ( .A(SITRAN_CMD1[9]), .B(n1642), .C(QTRAN_CMD1[9]), .D(n1617), 
        .E(ITRAN_CMD1[9]), .F(n1628), .Y(TRAN_CMD1[9]) );
    zao222b U157 ( .A(SITRAN_CMD1[10]), .B(n1643), .C(QTRAN_CMD1[10]), .D(
        n1648), .E(ITRAN_CMD1[10]), .F(n1635), .Y(TRAN_CMD1[10]) );
    zao222b U158 ( .A(SITRAN_CMD1[11]), .B(n1623), .C(QTRAN_CMD1[11]), .D(
        n1649), .E(ITRAN_CMD1[11]), .F(n1627), .Y(TRAN_CMD1[11]) );
    zao222b U159 ( .A(SITRAN_CMD1[12]), .B(n1623), .C(QTRAN_CMD1[12]), .D(
        n1617), .E(ITRAN_CMD1[12]), .F(n1635), .Y(TRAN_CMD1[12]) );
    zao222b U160 ( .A(SITRAN_CMD1[13]), .B(n1624), .C(QTRAN_CMD1[13]), .D(
        n1649), .E(ITRAN_CMD1[13]), .F(n1628), .Y(TRAN_CMD1[13]) );
    zao222b U161 ( .A(SITRAN_CMD1[14]), .B(n1623), .C(QTRAN_CMD1[14]), .D(
        n1617), .E(ITRAN_CMD1[14]), .F(n1628), .Y(TRAN_CMD1[14]) );
    zao222b U162 ( .A(SITRAN_CMD1[15]), .B(n1642), .C(QTRAN_CMD1[15]), .D(
        n1651), .E(ITRAN_CMD1[15]), .F(n1627), .Y(TRAN_CMD1[15]) );
    zao222b U163 ( .A(SITRAN_CMD1[16]), .B(n1612), .C(QTRAN_CMD1[16]), .D(
        n1648), .E(ITRAN_CMD1[16]), .F(n1637), .Y(TRAN_CMD1[16]) );
    zao222b U164 ( .A(SITRAN_CMD1[17]), .B(n1624), .C(QTRAN_CMD1[17]), .D(
        n1651), .E(ITRAN_CMD1[17]), .F(n1627), .Y(TRAN_CMD1[17]) );
    zao222b U165 ( .A(SITRAN_CMD1[18]), .B(n1641), .C(QTRAN_CMD1[18]), .D(
        n1617), .E(ITRAN_CMD1[18]), .F(n1637), .Y(TRAN_CMD1[18]) );
    zao222b U166 ( .A(SITRAN_CMD1[19]), .B(n1642), .C(QTRAN_CMD1[19]), .D(
        n1618), .E(ITRAN_CMD1[19]), .F(n1616), .Y(TRAN_CMD1[19]) );
    zao222b U167 ( .A(SITRAN_CMD1[20]), .B(n1642), .C(QTRAN_CMD1[20]), .D(
        n1618), .E(ITRAN_CMD1[20]), .F(n1616), .Y(TRAN_CMD1[20]) );
    zao222b U168 ( .A(SITRAN_CMD1[21]), .B(n1624), .C(QTRAN_CMD1[21]), .D(
        n1617), .E(ITRAN_CMD1[21]), .F(n1627), .Y(TRAN_CMD1[21]) );
    zao222b U169 ( .A(SITRAN_CMD1[22]), .B(n1643), .C(QTRAN_CMD1[22]), .D(
        n1618), .E(ITRAN_CMD1[22]), .F(n1616), .Y(TRAN_CMD1[22]) );
    zao222b U170 ( .A(SITRAN_CMD1[23]), .B(n1624), .C(QTRAN_CMD1[23]), .D(
        n1648), .E(ITRAN_CMD1[23]), .F(n1628), .Y(TRAN_CMD1[23]) );
    zao222b U171 ( .A(SITRAN_CMD1[24]), .B(n1643), .C(QTRAN_CMD1[24]), .D(
        n1651), .E(ITRAN_CMD1[24]), .F(n1636), .Y(TRAN_CMD1[24]) );
    zao222b U172 ( .A(SITRAN_CMD1[25]), .B(n1643), .C(QTRAN_CMD1[25]), .D(
        n1649), .E(ITRAN_CMD1[25]), .F(n1616), .Y(TRAN_CMD1[25]) );
    zao222b U173 ( .A(SITRAN_CMD1[26]), .B(n1643), .C(QTRAN_CMD1[26]), .D(
        n1650), .E(ITRAN_CMD1[26]), .F(n1627), .Y(TRAN_CMD1[26]) );
    zao222b U174 ( .A(SITRAN_CMD1[27]), .B(n1642), .C(QTRAN_CMD1[27]), .D(
        n1617), .E(ITRAN_CMD1[27]), .F(n1616), .Y(TRAN_CMD1[27]) );
    zao222b U175 ( .A(SITRAN_CMD1[28]), .B(n1612), .C(QTRAN_CMD1[28]), .D(
        n1648), .E(ITRAN_CMD1[28]), .F(n1635), .Y(TRAN_CMD1[28]) );
    zao222b U176 ( .A(SITRAN_CMD1[29]), .B(n1624), .C(QTRAN_CMD1[29]), .D(
        n1651), .E(ITRAN_CMD1[29]), .F(n1635), .Y(TRAN_CMD1[29]) );
    zao222b U177 ( .A(SITRAN_CMD1[30]), .B(n1642), .C(QTRAN_CMD1[30]), .D(
        n1651), .E(ITRAN_CMD1[30]), .F(n1616), .Y(TRAN_CMD1[30]) );
    zao222b U178 ( .A(SITRAN_CMD1[31]), .B(n1643), .C(QTRAN_CMD1[31]), .D(
        n1617), .E(ITRAN_CMD1[31]), .F(n1627), .Y(TRAN_CMD1[31]) );
    zao222b U179 ( .A(SITRAN_CMD1[32]), .B(n1623), .C(QTRAN_CMD1[32]), .D(
        n1650), .E(ITRAN_CMD1[32]), .F(n1635), .Y(TRAN_CMD1[32]) );
    zao222b U180 ( .A(SITRAN_CMD1[33]), .B(n1612), .C(QTRAN_CMD1[33]), .D(
        n1649), .E(ITRAN_CMD1[33]), .F(n1627), .Y(TRAN_CMD1[33]) );
    zao222b U181 ( .A(SITRAN_CMD1[34]), .B(n1624), .C(QTRAN_CMD1[34]), .D(
        n1648), .E(ITRAN_CMD1[34]), .F(n1616), .Y(TRAN_CMD1[34]) );
    zao222b U182 ( .A(SITRAN_CMD1[35]), .B(n1642), .C(QTRAN_CMD1[35]), .D(
        n1651), .E(ITRAN_CMD1[35]), .F(n1635), .Y(TRAN_CMD1[35]) );
    zao222b U183 ( .A(SITRAN_CMD1[36]), .B(n1624), .C(QTRAN_CMD1[36]), .D(
        n1651), .E(ITRAN_CMD1[36]), .F(n1637), .Y(TRAN_CMD1[36]) );
    zao222b U184 ( .A(SITRAN_CMD1[37]), .B(n1623), .C(QTRAN_CMD1[37]), .D(
        n1617), .E(ITRAN_CMD1[37]), .F(n1628), .Y(TRAN_CMD1[37]) );
    zao222b U185 ( .A(SITRAN_CMD1[38]), .B(n1623), .C(QTRAN_CMD1[38]), .D(
        n1650), .E(ITRAN_CMD1[38]), .F(n1627), .Y(TRAN_CMD1[38]) );
    zao222b U186 ( .A(SITRAN_CMD1[39]), .B(n1624), .C(QTRAN_CMD1[39]), .D(
        n1651), .E(ITRAN_CMD1[39]), .F(n1636), .Y(TRAN_CMD1[39]) );
    zao222b U187 ( .A(SITRAN_CMD1[40]), .B(n1624), .C(QTRAN_CMD1[40]), .D(
        n1648), .E(ITRAN_CMD1[40]), .F(n1628), .Y(TRAN_CMD1[40]) );
    zao222b U188 ( .A(SITRAN_CMD1[41]), .B(n1642), .C(QTRAN_CMD1[41]), .D(
        n1618), .E(ITRAN_CMD1[41]), .F(n1637), .Y(TRAN_CMD1[41]) );
    zao222b U189 ( .A(SITRAN_CMD1[42]), .B(n1641), .C(QTRAN_CMD1[42]), .D(
        n1617), .E(ITRAN_CMD1[42]), .F(n1616), .Y(TRAN_CMD1[42]) );
    zao222b U190 ( .A(SITRAN_CMD1[43]), .B(n1623), .C(QTRAN_CMD1[43]), .D(
        n1648), .E(ITRAN_CMD1[43]), .F(n1636), .Y(TRAN_CMD1[43]) );
    zao222b U191 ( .A(SITRAN_CMD1[44]), .B(n1642), .C(QTRAN_CMD1[44]), .D(
        n1649), .E(ITRAN_CMD1[44]), .F(n1636), .Y(TRAN_CMD1[44]) );
    zao222b U192 ( .A(SITRAN_CMD1[45]), .B(n1641), .C(QTRAN_CMD1[45]), .D(
        n1649), .E(ITRAN_CMD1[45]), .F(n1628), .Y(TRAN_CMD1[45]) );
    zao222b U193 ( .A(SITRAN_CMD1[46]), .B(n1642), .C(QTRAN_CMD1[46]), .D(
        n1618), .E(ITRAN_CMD1[46]), .F(n1627), .Y(TRAN_CMD1[46]) );
    zao222b U194 ( .A(SITRAN_CMD1[47]), .B(n1624), .C(QTRAN_CMD1[47]), .D(
        n1650), .E(ITRAN_CMD1[47]), .F(n1616), .Y(TRAN_CMD1[47]) );
    zao222b U195 ( .A(SITRAN_CMD1[48]), .B(n1641), .C(QTRAN_CMD1[48]), .D(
        n1650), .E(ITRAN_CMD1[48]), .F(n1637), .Y(TRAN_CMD1[48]) );
    zao222b U196 ( .A(SITRAN_CMD1[49]), .B(n1641), .C(QTRAN_CMD1[49]), .D(
        n1617), .E(ITRAN_CMD1[49]), .F(n1637), .Y(TRAN_CMD1[49]) );
    zao222b U197 ( .A(SITRAN_CMD1[50]), .B(n1624), .C(QTRAN_CMD1[50]), .D(
        n1650), .E(ITRAN_CMD1[50]), .F(n1628), .Y(TRAN_CMD1[50]) );
    zao222b U198 ( .A(SITRAN_CMD1[51]), .B(n1643), .C(QTRAN_CMD1[51]), .D(
        n1649), .E(ITRAN_CMD1[51]), .F(n1636), .Y(TRAN_CMD1[51]) );
    zao222b U199 ( .A(SITRAN_CMD1[52]), .B(n1643), .C(QTRAN_CMD1[52]), .D(
        n1651), .E(ITRAN_CMD1[52]), .F(n1628), .Y(TRAN_CMD1[52]) );
    zao222b U200 ( .A(SITRAN_CMD1[53]), .B(n1612), .C(QTRAN_CMD1[53]), .D(
        n1618), .E(ITRAN_CMD1[53]), .F(n1627), .Y(TRAN_CMD1[53]) );
    zao222b U201 ( .A(SITRAN_CMD1[54]), .B(n1641), .C(QTRAN_CMD1[54]), .D(
        n1650), .E(ITRAN_CMD1[54]), .F(n1635), .Y(TRAN_CMD1[54]) );
    zao222b U202 ( .A(SITRAN_CMD1[55]), .B(n1643), .C(QTRAN_CMD1[55]), .D(
        n1648), .E(ITRAN_CMD1[55]), .F(n1636), .Y(TRAN_CMD1[55]) );
    zao222b U203 ( .A(SITRAN_CMD1[56]), .B(n1642), .C(QTRAN_CMD1[56]), .D(
        n1617), .E(ITRAN_CMD1[56]), .F(n1636), .Y(TRAN_CMD1[56]) );
    zao222b U204 ( .A(SITRAN_CMD1[57]), .B(n1623), .C(QTRAN_CMD1[57]), .D(
        n1617), .E(ITRAN_CMD1[57]), .F(n1637), .Y(TRAN_CMD1[57]) );
    zao222b U205 ( .A(SITRAN_CMD1[58]), .B(n1623), .C(QTRAN_CMD1[58]), .D(
        n1650), .E(ITRAN_CMD1[58]), .F(n1616), .Y(TRAN_CMD1[58]) );
    zao222b U206 ( .A(SITRAN_CMD1[59]), .B(n1641), .C(QTRAN_CMD1[59]), .D(
        n1618), .E(ITRAN_CMD1[59]), .F(n1628), .Y(TRAN_CMD1[59]) );
    zao222b U207 ( .A(SITRAN_CMD1[60]), .B(n1612), .C(QTRAN_CMD1[60]), .D(
        n1648), .E(ITRAN_CMD1[60]), .F(n1616), .Y(TRAN_CMD1[60]) );
    zao222b U208 ( .A(SITRAN_CMD1[61]), .B(n1641), .C(QTRAN_CMD1[61]), .D(
        n1649), .E(ITRAN_CMD1[61]), .F(n1635), .Y(TRAN_CMD1[61]) );
    zao222b U209 ( .A(SITRAN_CMD1[62]), .B(n1624), .C(QTRAN_CMD1[62]), .D(
        n1650), .E(ITRAN_CMD1[62]), .F(n1616), .Y(TRAN_CMD1[62]) );
    zao222b U210 ( .A(SITRAN_CMD1[63]), .B(n1624), .C(QTRAN_CMD1[63]), .D(
        n1651), .E(ITRAN_CMD1[63]), .F(n1637), .Y(TRAN_CMD1[63]) );
    zao222b U211 ( .A(SITRAN_CMD1[64]), .B(n1641), .C(QTRAN_CMD1[64]), .D(
        n1650), .E(ITRAN_CMD1[64]), .F(n1616), .Y(TRAN_CMD1[64]) );
    zao222b U212 ( .A(SITRAN_CMD1[65]), .B(n1612), .C(QTRAN_CMD1[65]), .D(
        n1649), .E(ITRAN_CMD1[65]), .F(n1616), .Y(TRAN_CMD1[65]) );
    zao222b U213 ( .A(SITRAN_CMD1[66]), .B(n1643), .C(QTRAN_CMD1[66]), .D(
        n1648), .E(ITRAN_CMD1[66]), .F(n1637), .Y(TRAN_CMD1[66]) );
    zao222b U214 ( .A(SITRAN_CMD1[67]), .B(n1612), .C(QTRAN_CMD1[67]), .D(
        n1649), .E(ITRAN_CMD1[67]), .F(n1627), .Y(TRAN_CMD1[67]) );
    zao222b U215 ( .A(SITRAN_CMD1[68]), .B(n1642), .C(QTRAN_CMD1[68]), .D(
        n1648), .E(ITRAN_CMD1[68]), .F(n1636), .Y(TRAN_CMD1[68]) );
    zao222b U216 ( .A(SITRAN_CMD1[69]), .B(n1641), .C(QTRAN_CMD1[69]), .D(
        n1617), .E(ITRAN_CMD1[69]), .F(n1637), .Y(TRAN_CMD1[69]) );
    zao222b U217 ( .A(SITRAN_CMD1[70]), .B(n1623), .C(QTRAN_CMD1[70]), .D(
        n1648), .E(ITRAN_CMD1[70]), .F(n1627), .Y(TRAN_CMD1[70]) );
    zao222b U218 ( .A(SITRAN_CMD1[71]), .B(n1643), .C(QTRAN_CMD1[71]), .D(
        n1651), .E(ITRAN_CMD1[71]), .F(n1636), .Y(TRAN_CMD1[71]) );
    zao222b U219 ( .A(SITRAN_CMD1[72]), .B(n1643), .C(QTRAN_CMD1[72]), .D(
        n1648), .E(ITRAN_CMD1[72]), .F(n1628), .Y(TRAN_CMD1[72]) );
    zao222b U220 ( .A(SITRAN_CMD1[73]), .B(n1612), .C(QTRAN_CMD1[73]), .D(
        n1650), .E(ITRAN_CMD1[73]), .F(n1635), .Y(TRAN_CMD1[73]) );
    zao222b U221 ( .A(SITRAN_CMD1[74]), .B(n1642), .C(QTRAN_CMD1[74]), .D(
        n1650), .E(ITRAN_CMD1[74]), .F(n1628), .Y(TRAN_CMD1[74]) );
    zao222b U222 ( .A(SITRAN_CMD1[75]), .B(n1612), .C(QTRAN_CMD1[75]), .D(
        n1618), .E(ITRAN_CMD1[75]), .F(n1637), .Y(TRAN_CMD1[75]) );
    zao222b U223 ( .A(SITRAN_CMD1[76]), .B(n1612), .C(QTRAN_CMD1[76]), .D(
        n1651), .E(ITRAN_CMD1[76]), .F(n1616), .Y(TRAN_CMD1[76]) );
    zao222b U224 ( .A(SITRAN_CMD1[77]), .B(n1623), .C(QTRAN_CMD1[77]), .D(
        n1648), .E(ITRAN_CMD1[77]), .F(n1636), .Y(TRAN_CMD1[77]) );
    zao222b U225 ( .A(SITRAN_CMD1[78]), .B(n1642), .C(QTRAN_CMD1[78]), .D(
        n1618), .E(ITRAN_CMD1[78]), .F(n1627), .Y(TRAN_CMD1[78]) );
    zao222b U226 ( .A(SITRAN_CMD1[79]), .B(n1623), .C(QTRAN_CMD1[79]), .D(
        n1617), .E(ITRAN_CMD1[79]), .F(n1635), .Y(TRAN_CMD1[79]) );
    zao222b U227 ( .A(SITRAN_CMD1[80]), .B(n1641), .C(QTRAN_CMD1[80]), .D(
        n1649), .E(ITRAN_CMD1[80]), .F(n1637), .Y(TRAN_CMD1[80]) );
    zao222b U228 ( .A(SITRAN_CMD1[81]), .B(n1642), .C(QTRAN_CMD1[81]), .D(
        n1617), .E(ITRAN_CMD1[81]), .F(n1637), .Y(TRAN_CMD1[81]) );
    zao222b U229 ( .A(SITRAN_CMD1[82]), .B(n1624), .C(QTRAN_CMD1[82]), .D(
        n1618), .E(ITRAN_CMD1[82]), .F(n1636), .Y(TRAN_CMD1[82]) );
    zao222b U230 ( .A(SITRAN_CMD1[83]), .B(n1641), .C(QTRAN_CMD1[83]), .D(
        n1649), .E(ITRAN_CMD1[83]), .F(n1636), .Y(TRAN_CMD1[83]) );
    zao222b U231 ( .A(SITRAN_CMD1[84]), .B(n1612), .C(QTRAN_CMD1[84]), .D(
        n1650), .E(ITRAN_CMD1[84]), .F(n1616), .Y(TRAN_CMD1[84]) );
    zao222b U232 ( .A(SITRAN_CMD1[85]), .B(n1641), .C(QTRAN_CMD1[85]), .D(
        n1651), .E(ITRAN_CMD1[85]), .F(n1635), .Y(TRAN_CMD1[85]) );
    zao222b U233 ( .A(SITRAN_CMD1[86]), .B(n1623), .C(QTRAN_CMD1[86]), .D(
        n1649), .E(ITRAN_CMD1[86]), .F(n1616), .Y(TRAN_CMD1[86]) );
    zao222b U234 ( .A(SITRAN_CMD1[87]), .B(n1643), .C(QTRAN_CMD1[87]), .D(
        n1650), .E(ITRAN_CMD1[87]), .F(n1637), .Y(TRAN_CMD1[87]) );
    zao222b U235 ( .A(SITRAN_CMD1[88]), .B(n1612), .C(QTRAN_CMD1[88]), .D(
        n1651), .E(ITRAN_CMD1[88]), .F(n1628), .Y(TRAN_CMD1[88]) );
    zao222b U236 ( .A(SITRAN_CMD1[89]), .B(n1624), .C(QTRAN_CMD1[89]), .D(
        n1648), .E(ITRAN_CMD1[89]), .F(n1627), .Y(TRAN_CMD1[89]) );
    zao222b U237 ( .A(SITRAN_CMD1[90]), .B(n1643), .C(QTRAN_CMD1[90]), .D(
        n1649), .E(ITRAN_CMD1[90]), .F(n1627), .Y(TRAN_CMD1[90]) );
    zao222b U238 ( .A(SITRAN_CMD1[91]), .B(n1612), .C(QTRAN_CMD1[91]), .D(
        n1618), .E(ITRAN_CMD1[91]), .F(n1627), .Y(TRAN_CMD1[91]) );
    zao222b U239 ( .A(SITRAN_CMD1[92]), .B(n1623), .C(QTRAN_CMD1[92]), .D(
        n1651), .E(ITRAN_CMD1[92]), .F(n1637), .Y(TRAN_CMD1[92]) );
    zao222b U240 ( .A(SITRAN_CMD1[93]), .B(n1612), .C(QTRAN_CMD1[93]), .D(
        n1651), .E(ITRAN_CMD1[93]), .F(n1636), .Y(TRAN_CMD1[93]) );
    zao222b U241 ( .A(SITRAN_CMD1[94]), .B(n1624), .C(QTRAN_CMD1[94]), .D(
        n1618), .E(ITRAN_CMD1[94]), .F(n1636), .Y(TRAN_CMD1[94]) );
    zao222b U242 ( .A(SITRAN_CMD1[95]), .B(n1642), .C(QTRAN_CMD1[95]), .D(
        n1650), .E(ITRAN_CMD1[95]), .F(n1628), .Y(TRAN_CMD1[95]) );
    zao222b U243 ( .A(SITRAN_CMD1[96]), .B(n1641), .C(QTRAN_CMD1[96]), .D(
        n1650), .E(ITRAN_CMD1[96]), .F(n1635), .Y(TRAN_CMD1[96]) );
    zao222b U244 ( .A(SITRAN_CMD1[97]), .B(n1623), .C(QTRAN_CMD1[97]), .D(
        n1617), .E(ITRAN_CMD1[97]), .F(n1627), .Y(TRAN_CMD1[97]) );
    zao222b U245 ( .A(SITRAN_CMD1[98]), .B(n1643), .C(QTRAN_CMD1[98]), .D(
        n1618), .E(ITRAN_CMD1[98]), .F(n1637), .Y(TRAN_CMD1[98]) );
    zao222b U246 ( .A(n1624), .B(SITRAN_CMD1[99]), .C(n1618), .D(QTRAN_CMD1
        [99]), .E(n1616), .F(ITRAN_CMD1[99]), .Y(TRAN_CMD1[99]) );
    zao222b U247 ( .A(SITRAN_CMD1[100]), .B(n1643), .C(QTRAN_CMD1[100]), .D(
        n1617), .E(ITRAN_CMD1[100]), .F(n1635), .Y(TRAN_CMD1[100]) );
    zao222b U248 ( .A(SITRAN_CMD1[101]), .B(n1642), .C(QTRAN_CMD1[101]), .D(
        n1617), .E(ITRAN_CMD1[101]), .F(n1628), .Y(TRAN_CMD1[101]) );
    zao222b U249 ( .A(SITRAN_CMD1[102]), .B(n1623), .C(QTRAN_CMD1[102]), .D(
        n1649), .E(ITRAN_CMD1[102]), .F(n1636), .Y(TRAN_CMD1[102]) );
    zao222b U250 ( .A(SITRAN_CMD1[103]), .B(n1612), .C(QTRAN_CMD1[103]), .D(
        n1618), .E(ITRAN_CMD1[103]), .F(n1635), .Y(TRAN_CMD1[103]) );
    zao222b U251 ( .A(SITRAN_CMD1[104]), .B(n1641), .C(QTRAN_CMD1[104]), .D(
        n1617), .E(ITRAN_CMD1[104]), .F(n1628), .Y(TRAN_CMD1[104]) );
    zan2b U252 ( .A(CRCERR), .B(n1629), .Y(CRCERR2) );
    zan2b U253 ( .A(BABBLE), .B(n1629), .Y(BABBLE2) );
    zan2b U254 ( .A(PIDERR), .B(n1629), .Y(PIDERR2) );
    zan2b U255 ( .A(TMOUT), .B(n1629), .Y(TMOUT2) );
    zan2b U256 ( .A(n1629), .B(TOGMATCH), .Y(TOGMATCH2) );
    zan2b U257 ( .A(RXNAK), .B(n1629), .Y(RXNAK2) );
    zan2b U258 ( .A(RXNYET), .B(USBDMA_SEL[1]), .Y(RXNYET2) );
    zan2b U259 ( .A(RXSTALL), .B(USBDMA_SEL[1]), .Y(RXSTALL2) );
    zan2b U260 ( .A(RXACK), .B(USBDMA_SEL[1]), .Y(RXACK2) );
    zan2b U261 ( .A(RXDATA0), .B(USBDMA_SEL[1]), .Y(RXDATA02) );
    zan2b U262 ( .A(RXDATA1), .B(n1629), .Y(RXDATA12) );
    zan2b U263 ( .A(RXDATA2), .B(n1629), .Y(RXDATA22) );
    zan2b U264 ( .A(RXMDATA), .B(USBDMA_SEL[1]), .Y(RXMDATA2) );
    zan2b U265 ( .A(RXPIDERR), .B(n1629), .Y(RXPIDERR2) );
    zan2b U266 ( .A(SPD), .B(n1629), .Y(SPD2) );
    zan2b U267 ( .A(ACTLEN[10]), .B(USBDMA_SEL[1]), .Y(ACTLEN2[10]) );
    zan2b U268 ( .A(ACTLEN[9]), .B(n1629), .Y(ACTLEN2[9]) );
    zan2b U269 ( .A(ACTLEN[8]), .B(USBDMA_SEL[1]), .Y(ACTLEN2[8]) );
    zan2b U270 ( .A(ACTLEN[7]), .B(USBDMA_SEL[1]), .Y(ACTLEN2[7]) );
    zan2b U271 ( .A(ACTLEN[6]), .B(n1629), .Y(ACTLEN2[6]) );
    zan2b U272 ( .A(ACTLEN[5]), .B(n1629), .Y(ACTLEN2[5]) );
    zan2b U273 ( .A(ACTLEN[4]), .B(n1629), .Y(ACTLEN2[4]) );
    zan2b U274 ( .A(ACTLEN[3]), .B(n1629), .Y(ACTLEN2[3]) );
    zan2b U275 ( .A(ACTLEN[2]), .B(n1629), .Y(ACTLEN2[2]) );
    zan2b U276 ( .A(ACTLEN[1]), .B(n1629), .Y(ACTLEN2[1]) );
    zan2b U277 ( .A(ACTLEN[0]), .B(n1629), .Y(ACTLEN2[0]) );
    zao222b U278 ( .A(SITRAN_CMD2[0]), .B(n1620), .C(QTRAN_CMD2[0]), .D(n1654), 
        .E(ITRAN_CMD2[0]), .F(n1639), .Y(TRAN_CMD2[0]) );
    zao222b U279 ( .A(SITRAN_CMD2[1]), .B(n1620), .C(QTRAN_CMD2[1]), .D(n1656), 
        .E(ITRAN_CMD2[1]), .F(n1640), .Y(TRAN_CMD2[1]) );
    zao222b U280 ( .A(SITRAN_CMD2[2]), .B(n1644), .C(QTRAN_CMD2[2]), .D(n1655), 
        .E(ITRAN_CMD2[2]), .F(n1639), .Y(TRAN_CMD2[2]) );
    zao222b U281 ( .A(SITRAN_CMD2[3]), .B(n1619), .C(QTRAN_CMD2[3]), .D(n1622), 
        .E(ITRAN_CMD2[3]), .F(n1639), .Y(TRAN_CMD2[3]) );
    zao222b U282 ( .A(SITRAN_CMD2[4]), .B(n1646), .C(QTRAN_CMD2[4]), .D(n1654), 
        .E(ITRAN_CMD2[4]), .F(n1614), .Y(TRAN_CMD2[4]) );
    zao222b U283 ( .A(SITRAN_CMD2[5]), .B(n1619), .C(QTRAN_CMD2[5]), .D(n1622), 
        .E(ITRAN_CMD2[5]), .F(n1625), .Y(TRAN_CMD2[5]) );
    zao222b U284 ( .A(SITRAN_CMD2[6]), .B(n1610), .C(QTRAN_CMD2[6]), .D(n1656), 
        .E(ITRAN_CMD2[6]), .F(n1614), .Y(TRAN_CMD2[6]) );
    zao222b U285 ( .A(SITRAN_CMD2[7]), .B(n1645), .C(QTRAN_CMD2[7]), .D(n1653), 
        .E(ITRAN_CMD2[7]), .F(n1640), .Y(TRAN_CMD2[7]) );
    zao222b U286 ( .A(SITRAN_CMD2[8]), .B(n1644), .C(QTRAN_CMD2[8]), .D(n1656), 
        .E(ITRAN_CMD2[8]), .F(n1626), .Y(TRAN_CMD2[8]) );
    zao222b U287 ( .A(SITRAN_CMD2[9]), .B(n1645), .C(QTRAN_CMD2[9]), .D(n1621), 
        .E(ITRAN_CMD2[9]), .F(n1638), .Y(TRAN_CMD2[9]) );
    zao222b U288 ( .A(SITRAN_CMD2[10]), .B(n1646), .C(QTRAN_CMD2[10]), .D(
        n1653), .E(ITRAN_CMD2[10]), .F(n1614), .Y(TRAN_CMD2[10]) );
    zao222b U289 ( .A(SITRAN_CMD2[11]), .B(n1619), .C(QTRAN_CMD2[11]), .D(
        n1654), .E(ITRAN_CMD2[11]), .F(n1614), .Y(TRAN_CMD2[11]) );
    zao222b U290 ( .A(SITRAN_CMD2[12]), .B(n1619), .C(QTRAN_CMD2[12]), .D(
        n1621), .E(ITRAN_CMD2[12]), .F(n1640), .Y(TRAN_CMD2[12]) );
    zao222b U291 ( .A(SITRAN_CMD2[13]), .B(n1620), .C(QTRAN_CMD2[13]), .D(
        n1654), .E(ITRAN_CMD2[13]), .F(n1626), .Y(TRAN_CMD2[13]) );
    zao222b U292 ( .A(SITRAN_CMD2[14]), .B(n1619), .C(QTRAN_CMD2[14]), .D(
        n1621), .E(ITRAN_CMD2[14]), .F(n1640), .Y(TRAN_CMD2[14]) );
    zao222b U293 ( .A(SITRAN_CMD2[15]), .B(n1645), .C(QTRAN_CMD2[15]), .D(
        n1656), .E(ITRAN_CMD2[15]), .F(n1639), .Y(TRAN_CMD2[15]) );
    zao222b U294 ( .A(SITRAN_CMD2[16]), .B(n1610), .C(QTRAN_CMD2[16]), .D(
        n1653), .E(ITRAN_CMD2[16]), .F(n1638), .Y(TRAN_CMD2[16]) );
    zao222b U295 ( .A(SITRAN_CMD2[17]), .B(n1620), .C(QTRAN_CMD2[17]), .D(
        n1656), .E(ITRAN_CMD2[17]), .F(n1625), .Y(TRAN_CMD2[17]) );
    zao222b U296 ( .A(SITRAN_CMD2[18]), .B(n1644), .C(QTRAN_CMD2[18]), .D(
        n1621), .E(ITRAN_CMD2[18]), .F(n1639), .Y(TRAN_CMD2[18]) );
    zao222b U297 ( .A(SITRAN_CMD2[19]), .B(n1645), .C(QTRAN_CMD2[19]), .D(
        n1622), .E(ITRAN_CMD2[19]), .F(n1625), .Y(TRAN_CMD2[19]) );
    zao222b U298 ( .A(SITRAN_CMD2[20]), .B(n1645), .C(QTRAN_CMD2[20]), .D(
        n1622), .E(ITRAN_CMD2[20]), .F(n1638), .Y(TRAN_CMD2[20]) );
    zao222b U299 ( .A(SITRAN_CMD2[21]), .B(n1620), .C(QTRAN_CMD2[21]), .D(
        n1621), .E(ITRAN_CMD2[21]), .F(n1638), .Y(TRAN_CMD2[21]) );
    zao222b U300 ( .A(SITRAN_CMD2[22]), .B(n1646), .C(QTRAN_CMD2[22]), .D(
        n1622), .E(ITRAN_CMD2[22]), .F(n1626), .Y(TRAN_CMD2[22]) );
    zao222b U301 ( .A(SITRAN_CMD2[23]), .B(n1620), .C(QTRAN_CMD2[23]), .D(
        n1653), .E(ITRAN_CMD2[23]), .F(n1614), .Y(TRAN_CMD2[23]) );
    zao222b U302 ( .A(SITRAN_CMD2[24]), .B(n1646), .C(QTRAN_CMD2[24]), .D(
        n1656), .E(ITRAN_CMD2[24]), .F(n1626), .Y(TRAN_CMD2[24]) );
    zao222b U303 ( .A(SITRAN_CMD2[25]), .B(n1646), .C(QTRAN_CMD2[25]), .D(
        n1654), .E(ITRAN_CMD2[25]), .F(n1640), .Y(TRAN_CMD2[25]) );
    zao222b U304 ( .A(SITRAN_CMD2[26]), .B(n1646), .C(QTRAN_CMD2[26]), .D(
        n1655), .E(ITRAN_CMD2[26]), .F(n1614), .Y(TRAN_CMD2[26]) );
    zao222b U305 ( .A(SITRAN_CMD2[27]), .B(n1645), .C(QTRAN_CMD2[27]), .D(
        n1621), .E(ITRAN_CMD2[27]), .F(n1625), .Y(TRAN_CMD2[27]) );
    zao222b U306 ( .A(SITRAN_CMD2[28]), .B(n1610), .C(QTRAN_CMD2[28]), .D(
        n1653), .E(ITRAN_CMD2[28]), .F(n1625), .Y(TRAN_CMD2[28]) );
    zao222b U307 ( .A(SITRAN_CMD2[29]), .B(n1620), .C(QTRAN_CMD2[29]), .D(
        n1656), .E(ITRAN_CMD2[29]), .F(n1638), .Y(TRAN_CMD2[29]) );
    zao222b U308 ( .A(SITRAN_CMD2[30]), .B(n1645), .C(QTRAN_CMD2[30]), .D(
        n1656), .E(ITRAN_CMD2[30]), .F(n1626), .Y(TRAN_CMD2[30]) );
    zao222b U309 ( .A(SITRAN_CMD2[31]), .B(n1646), .C(QTRAN_CMD2[31]), .D(
        n1621), .E(ITRAN_CMD2[31]), .F(n1626), .Y(TRAN_CMD2[31]) );
    zao222b U310 ( .A(SITRAN_CMD2[32]), .B(n1619), .C(QTRAN_CMD2[32]), .D(
        n1655), .E(ITRAN_CMD2[32]), .F(n1640), .Y(TRAN_CMD2[32]) );
    zao222b U311 ( .A(SITRAN_CMD2[33]), .B(n1610), .C(QTRAN_CMD2[33]), .D(
        n1654), .E(ITRAN_CMD2[33]), .F(n1640), .Y(TRAN_CMD2[33]) );
    zao222b U312 ( .A(SITRAN_CMD2[34]), .B(n1620), .C(QTRAN_CMD2[34]), .D(
        n1653), .E(ITRAN_CMD2[34]), .F(n1614), .Y(TRAN_CMD2[34]) );
    zao222b U313 ( .A(SITRAN_CMD2[35]), .B(n1645), .C(QTRAN_CMD2[35]), .D(
        n1656), .E(ITRAN_CMD2[35]), .F(n1638), .Y(TRAN_CMD2[35]) );
    zao222b U314 ( .A(SITRAN_CMD2[36]), .B(n1620), .C(QTRAN_CMD2[36]), .D(
        n1656), .E(ITRAN_CMD2[36]), .F(n1638), .Y(TRAN_CMD2[36]) );
    zao222b U315 ( .A(SITRAN_CMD2[37]), .B(n1619), .C(QTRAN_CMD2[37]), .D(
        n1621), .E(ITRAN_CMD2[37]), .F(n1626), .Y(TRAN_CMD2[37]) );
    zao222b U316 ( .A(SITRAN_CMD2[38]), .B(n1619), .C(QTRAN_CMD2[38]), .D(
        n1655), .E(ITRAN_CMD2[38]), .F(n1640), .Y(TRAN_CMD2[38]) );
    zao222b U317 ( .A(SITRAN_CMD2[39]), .B(n1620), .C(QTRAN_CMD2[39]), .D(
        n1656), .E(ITRAN_CMD2[39]), .F(n1626), .Y(TRAN_CMD2[39]) );
    zao222b U318 ( .A(SITRAN_CMD2[40]), .B(n1620), .C(QTRAN_CMD2[40]), .D(
        n1653), .E(ITRAN_CMD2[40]), .F(n1640), .Y(TRAN_CMD2[40]) );
    zao222b U319 ( .A(SITRAN_CMD2[41]), .B(n1645), .C(QTRAN_CMD2[41]), .D(
        n1622), .E(ITRAN_CMD2[41]), .F(n1638), .Y(TRAN_CMD2[41]) );
    zao222b U320 ( .A(SITRAN_CMD2[42]), .B(n1644), .C(QTRAN_CMD2[42]), .D(
        n1621), .E(ITRAN_CMD2[42]), .F(n1640), .Y(TRAN_CMD2[42]) );
    zao222b U321 ( .A(SITRAN_CMD2[43]), .B(n1619), .C(QTRAN_CMD2[43]), .D(
        n1653), .E(ITRAN_CMD2[43]), .F(n1626), .Y(TRAN_CMD2[43]) );
    zao222b U322 ( .A(SITRAN_CMD2[44]), .B(n1645), .C(QTRAN_CMD2[44]), .D(
        n1654), .E(ITRAN_CMD2[44]), .F(n1639), .Y(TRAN_CMD2[44]) );
    zao222b U323 ( .A(SITRAN_CMD2[45]), .B(n1644), .C(QTRAN_CMD2[45]), .D(
        n1654), .E(ITRAN_CMD2[45]), .F(n1614), .Y(TRAN_CMD2[45]) );
    zao222b U324 ( .A(SITRAN_CMD2[46]), .B(n1645), .C(QTRAN_CMD2[46]), .D(
        n1622), .E(ITRAN_CMD2[46]), .F(n1625), .Y(TRAN_CMD2[46]) );
    zao222b U325 ( .A(SITRAN_CMD2[47]), .B(n1620), .C(QTRAN_CMD2[47]), .D(
        n1655), .E(ITRAN_CMD2[47]), .F(n1625), .Y(TRAN_CMD2[47]) );
    zao222b U326 ( .A(SITRAN_CMD2[48]), .B(n1644), .C(QTRAN_CMD2[48]), .D(
        n1655), .E(ITRAN_CMD2[48]), .F(n1638), .Y(TRAN_CMD2[48]) );
    zao222b U327 ( .A(SITRAN_CMD2[49]), .B(n1644), .C(QTRAN_CMD2[49]), .D(
        n1621), .E(ITRAN_CMD2[49]), .F(n1638), .Y(TRAN_CMD2[49]) );
    zao222b U328 ( .A(SITRAN_CMD2[50]), .B(n1620), .C(QTRAN_CMD2[50]), .D(
        n1655), .E(ITRAN_CMD2[50]), .F(n1626), .Y(TRAN_CMD2[50]) );
    zao222b U329 ( .A(SITRAN_CMD2[51]), .B(n1646), .C(QTRAN_CMD2[51]), .D(
        n1654), .E(ITRAN_CMD2[51]), .F(n1614), .Y(TRAN_CMD2[51]) );
    zao222b U330 ( .A(SITRAN_CMD2[52]), .B(n1646), .C(QTRAN_CMD2[52]), .D(
        n1656), .E(ITRAN_CMD2[52]), .F(n1626), .Y(TRAN_CMD2[52]) );
    zao222b U331 ( .A(SITRAN_CMD2[53]), .B(n1610), .C(QTRAN_CMD2[53]), .D(
        n1622), .E(ITRAN_CMD2[53]), .F(n1640), .Y(TRAN_CMD2[53]) );
    zao222b U332 ( .A(SITRAN_CMD2[54]), .B(n1644), .C(QTRAN_CMD2[54]), .D(
        n1655), .E(ITRAN_CMD2[54]), .F(n1639), .Y(TRAN_CMD2[54]) );
    zao222b U333 ( .A(SITRAN_CMD2[55]), .B(n1646), .C(QTRAN_CMD2[55]), .D(
        n1653), .E(ITRAN_CMD2[55]), .F(n1639), .Y(TRAN_CMD2[55]) );
    zao222b U334 ( .A(SITRAN_CMD2[56]), .B(n1645), .C(QTRAN_CMD2[56]), .D(
        n1621), .E(ITRAN_CMD2[56]), .F(n1626), .Y(TRAN_CMD2[56]) );
    zao222b U335 ( .A(SITRAN_CMD2[57]), .B(n1619), .C(QTRAN_CMD2[57]), .D(
        n1621), .E(ITRAN_CMD2[57]), .F(n1638), .Y(TRAN_CMD2[57]) );
    zao222b U336 ( .A(SITRAN_CMD2[58]), .B(n1619), .C(QTRAN_CMD2[58]), .D(
        n1655), .E(ITRAN_CMD2[58]), .F(n1639), .Y(TRAN_CMD2[58]) );
    zao222b U337 ( .A(SITRAN_CMD2[59]), .B(n1644), .C(QTRAN_CMD2[59]), .D(
        n1622), .E(ITRAN_CMD2[59]), .F(n1625), .Y(TRAN_CMD2[59]) );
    zao222b U338 ( .A(SITRAN_CMD2[60]), .B(n1610), .C(QTRAN_CMD2[60]), .D(
        n1653), .E(ITRAN_CMD2[60]), .F(n1639), .Y(TRAN_CMD2[60]) );
    zao222b U339 ( .A(SITRAN_CMD2[61]), .B(n1644), .C(QTRAN_CMD2[61]), .D(
        n1654), .E(ITRAN_CMD2[61]), .F(n1640), .Y(TRAN_CMD2[61]) );
    zao222b U340 ( .A(SITRAN_CMD2[62]), .B(n1620), .C(QTRAN_CMD2[62]), .D(
        n1655), .E(ITRAN_CMD2[62]), .F(n1625), .Y(TRAN_CMD2[62]) );
    zao222b U341 ( .A(SITRAN_CMD2[63]), .B(n1620), .C(QTRAN_CMD2[63]), .D(
        n1656), .E(ITRAN_CMD2[63]), .F(n1638), .Y(TRAN_CMD2[63]) );
    zao222b U342 ( .A(SITRAN_CMD2[64]), .B(n1644), .C(QTRAN_CMD2[64]), .D(
        n1655), .E(ITRAN_CMD2[64]), .F(n1640), .Y(TRAN_CMD2[64]) );
    zao222b U343 ( .A(SITRAN_CMD2[65]), .B(n1610), .C(QTRAN_CMD2[65]), .D(
        n1654), .E(ITRAN_CMD2[65]), .F(n1640), .Y(TRAN_CMD2[65]) );
    zao222b U344 ( .A(SITRAN_CMD2[66]), .B(n1646), .C(QTRAN_CMD2[66]), .D(
        n1653), .E(ITRAN_CMD2[66]), .F(n1625), .Y(TRAN_CMD2[66]) );
    zao222b U345 ( .A(SITRAN_CMD2[67]), .B(n1610), .C(QTRAN_CMD2[67]), .D(
        n1654), .E(ITRAN_CMD2[67]), .F(n1625), .Y(TRAN_CMD2[67]) );
    zao222b U346 ( .A(SITRAN_CMD2[68]), .B(n1645), .C(QTRAN_CMD2[68]), .D(
        n1653), .E(ITRAN_CMD2[68]), .F(n1614), .Y(TRAN_CMD2[68]) );
    zao222b U347 ( .A(SITRAN_CMD2[69]), .B(n1644), .C(QTRAN_CMD2[69]), .D(
        n1621), .E(ITRAN_CMD2[69]), .F(n1638), .Y(TRAN_CMD2[69]) );
    zao222b U348 ( .A(SITRAN_CMD2[70]), .B(n1619), .C(QTRAN_CMD2[70]), .D(
        n1653), .E(ITRAN_CMD2[70]), .F(n1614), .Y(TRAN_CMD2[70]) );
    zao222b U349 ( .A(SITRAN_CMD2[71]), .B(n1646), .C(QTRAN_CMD2[71]), .D(
        n1656), .E(ITRAN_CMD2[71]), .F(n1626), .Y(TRAN_CMD2[71]) );
    zao222b U350 ( .A(SITRAN_CMD2[72]), .B(n1646), .C(QTRAN_CMD2[72]), .D(
        n1653), .E(ITRAN_CMD2[72]), .F(n1614), .Y(TRAN_CMD2[72]) );
    zao222b U351 ( .A(SITRAN_CMD2[73]), .B(n1610), .C(QTRAN_CMD2[73]), .D(
        n1655), .E(ITRAN_CMD2[73]), .F(n1640), .Y(TRAN_CMD2[73]) );
    zao222b U352 ( .A(SITRAN_CMD2[74]), .B(n1645), .C(QTRAN_CMD2[74]), .D(
        n1655), .E(ITRAN_CMD2[74]), .F(n1639), .Y(TRAN_CMD2[74]) );
    zao222b U353 ( .A(SITRAN_CMD2[75]), .B(n1610), .C(QTRAN_CMD2[75]), .D(
        n1622), .E(ITRAN_CMD2[75]), .F(n1638), .Y(TRAN_CMD2[75]) );
    zao222b U354 ( .A(SITRAN_CMD2[76]), .B(n1610), .C(QTRAN_CMD2[76]), .D(
        n1656), .E(ITRAN_CMD2[76]), .F(n1625), .Y(TRAN_CMD2[76]) );
    zao222b U355 ( .A(SITRAN_CMD2[77]), .B(n1619), .C(QTRAN_CMD2[77]), .D(
        n1653), .E(ITRAN_CMD2[77]), .F(n1614), .Y(TRAN_CMD2[77]) );
    zao222b U356 ( .A(SITRAN_CMD2[78]), .B(n1645), .C(QTRAN_CMD2[78]), .D(
        n1622), .E(ITRAN_CMD2[78]), .F(n1639), .Y(TRAN_CMD2[78]) );
    zao222b U357 ( .A(SITRAN_CMD2[79]), .B(n1619), .C(QTRAN_CMD2[79]), .D(
        n1621), .E(ITRAN_CMD2[79]), .F(n1625), .Y(TRAN_CMD2[79]) );
    zao222b U358 ( .A(SITRAN_CMD2[80]), .B(n1644), .C(QTRAN_CMD2[80]), .D(
        n1654), .E(ITRAN_CMD2[80]), .F(n1614), .Y(TRAN_CMD2[80]) );
    zao222b U359 ( .A(SITRAN_CMD2[81]), .B(n1645), .C(QTRAN_CMD2[81]), .D(
        n1621), .E(ITRAN_CMD2[81]), .F(n1638), .Y(TRAN_CMD2[81]) );
    zao222b U360 ( .A(SITRAN_CMD2[82]), .B(n1620), .C(QTRAN_CMD2[82]), .D(
        n1622), .E(ITRAN_CMD2[82]), .F(n1626), .Y(TRAN_CMD2[82]) );
    zao222b U361 ( .A(SITRAN_CMD2[83]), .B(n1644), .C(QTRAN_CMD2[83]), .D(
        n1654), .E(ITRAN_CMD2[83]), .F(n1614), .Y(TRAN_CMD2[83]) );
    zao222b U362 ( .A(SITRAN_CMD2[84]), .B(n1610), .C(QTRAN_CMD2[84]), .D(
        n1655), .E(ITRAN_CMD2[84]), .F(n1639), .Y(TRAN_CMD2[84]) );
    zao222b U363 ( .A(SITRAN_CMD2[85]), .B(n1644), .C(QTRAN_CMD2[85]), .D(
        n1656), .E(ITRAN_CMD2[85]), .F(n1625), .Y(TRAN_CMD2[85]) );
    zao222b U364 ( .A(SITRAN_CMD2[86]), .B(n1619), .C(QTRAN_CMD2[86]), .D(
        n1654), .E(ITRAN_CMD2[86]), .F(n1626), .Y(TRAN_CMD2[86]) );
    zao222b U365 ( .A(SITRAN_CMD2[87]), .B(n1646), .C(QTRAN_CMD2[87]), .D(
        n1655), .E(ITRAN_CMD2[87]), .F(n1638), .Y(TRAN_CMD2[87]) );
    zao222b U366 ( .A(SITRAN_CMD2[88]), .B(n1610), .C(QTRAN_CMD2[88]), .D(
        n1656), .E(ITRAN_CMD2[88]), .F(n1640), .Y(TRAN_CMD2[88]) );
    zao222b U367 ( .A(SITRAN_CMD2[89]), .B(n1620), .C(QTRAN_CMD2[89]), .D(
        n1653), .E(ITRAN_CMD2[89]), .F(n1625), .Y(TRAN_CMD2[89]) );
    zao222b U368 ( .A(SITRAN_CMD2[90]), .B(n1646), .C(QTRAN_CMD2[90]), .D(
        n1654), .E(ITRAN_CMD2[90]), .F(n1625), .Y(TRAN_CMD2[90]) );
    zao222b U369 ( .A(SITRAN_CMD2[91]), .B(n1610), .C(QTRAN_CMD2[91]), .D(
        n1622), .E(ITRAN_CMD2[91]), .F(n1625), .Y(TRAN_CMD2[91]) );
    zao222b U370 ( .A(SITRAN_CMD2[92]), .B(n1619), .C(QTRAN_CMD2[92]), .D(
        n1656), .E(ITRAN_CMD2[92]), .F(n1638), .Y(TRAN_CMD2[92]) );
    zao222b U371 ( .A(SITRAN_CMD2[93]), .B(n1610), .C(QTRAN_CMD2[93]), .D(
        n1656), .E(ITRAN_CMD2[93]), .F(n1640), .Y(TRAN_CMD2[93]) );
    zao222b U372 ( .A(SITRAN_CMD2[94]), .B(n1620), .C(QTRAN_CMD2[94]), .D(
        n1622), .E(ITRAN_CMD2[94]), .F(n1614), .Y(TRAN_CMD2[94]) );
    zao222b U373 ( .A(SITRAN_CMD2[95]), .B(n1645), .C(QTRAN_CMD2[95]), .D(
        n1655), .E(ITRAN_CMD2[95]), .F(n1614), .Y(TRAN_CMD2[95]) );
    zao222b U374 ( .A(SITRAN_CMD2[96]), .B(n1644), .C(QTRAN_CMD2[96]), .D(
        n1655), .E(ITRAN_CMD2[96]), .F(n1625), .Y(TRAN_CMD2[96]) );
    zao222b U375 ( .A(SITRAN_CMD2[97]), .B(n1619), .C(QTRAN_CMD2[97]), .D(
        n1621), .E(ITRAN_CMD2[97]), .F(n1639), .Y(TRAN_CMD2[97]) );
    zao222b U376 ( .A(SITRAN_CMD2[98]), .B(n1646), .C(QTRAN_CMD2[98]), .D(
        n1622), .E(ITRAN_CMD2[98]), .F(n1638), .Y(TRAN_CMD2[98]) );
    zao222b U377 ( .A(n1620), .B(SITRAN_CMD2[99]), .C(n1622), .D(QTRAN_CMD2
        [99]), .E(n1640), .F(ITRAN_CMD2[99]), .Y(TRAN_CMD2[99]) );
    zao222b U378 ( .A(SITRAN_CMD2[100]), .B(n1646), .C(QTRAN_CMD2[100]), .D(
        n1621), .E(ITRAN_CMD2[100]), .F(n1614), .Y(TRAN_CMD2[100]) );
    zao222b U379 ( .A(SITRAN_CMD2[101]), .B(n1645), .C(QTRAN_CMD2[101]), .D(
        n1621), .E(ITRAN_CMD2[101]), .F(n1614), .Y(TRAN_CMD2[101]) );
    zao222b U380 ( .A(SITRAN_CMD2[102]), .B(n1619), .C(QTRAN_CMD2[102]), .D(
        n1654), .E(ITRAN_CMD2[102]), .F(n1626), .Y(TRAN_CMD2[102]) );
    zao222b U381 ( .A(SITRAN_CMD2[103]), .B(n1610), .C(QTRAN_CMD2[103]), .D(
        n1622), .E(ITRAN_CMD2[103]), .F(n1625), .Y(TRAN_CMD2[103]) );
    zao222b U382 ( .A(SITRAN_CMD2[104]), .B(n1644), .C(QTRAN_CMD2[104]), .D(
        n1621), .E(ITRAN_CMD2[104]), .F(n1639), .Y(TRAN_CMD2[104]) );
    zan2b U383 ( .A(PER_CMDSTART1), .B(n1633), .Y(QCMDSTART1) );
    zor3b U384 ( .A(SITDPARSING1), .B(ITDPARSING1), .C(QHPARSING1), .Y(
        TDPARSING1) );
    zan2b U385 ( .A(SITD_ACT2), .B(EHCI_MAC_EOT), .Y(SITD_MAC_EOT2) );
    zor3b U386 ( .A(SIBUI_GO1), .B(IBUI_GO1), .C(QBUI_GO1), .Y(BUI_GO1) );
    zor3b U387 ( .A(SIRXERR2), .B(IRXERR2), .C(QRXERR2), .Y(RXERR2) );
    zor3b U388 ( .A(SICMDSTART_REQ2), .B(ICMDSTART_REQ2), .C(QCMDSTART_REQ2), 
        .Y(PER_CMDSTART_REQ2) );
    zan2b U389 ( .A(n1679), .B(n1638), .Y(IPCIEND2) );
    zan2b U390 ( .A(TD_PARSE_GO1), .B(n1633), .Y(QH_PARSE_GO1) );
    zan2b U391 ( .A(EHCI_MAC_EOT), .B(QH_ACT2), .Y(QH_MAC_EOT2) );
    zan2b U392 ( .A(PER_CMDSTART2), .B(n1614), .Y(ICMDSTART2) );
    zor3b U393 ( .A(SICACHE_INVALID2), .B(ICACHE_INVALID2), .C(QCACHE_INVALID2
        ), .Y(CACHE_INVALID2) );
    zor3b U394 ( .A(SIHCIREQ2), .B(IHCIREQ2), .C(QHCIREQ2), .Y(TDHCIREQ2) );
    zor3b U395 ( .A(SIRXERR1), .B(IRXERR1), .C(QRXERR1), .Y(RXERR1) );
    zan2b U396 ( .A(TD_PARSE_GO2), .B(n1631), .Y(QH_PARSE_GO2) );
    zan2b U397 ( .A(EHCI_MAC_EOT), .B(QH_ACT1), .Y(QH_MAC_EOT1) );
    zor3b U398 ( .A(PARSEITDEND2), .B(PARSEQHEND2), .C(PARSESITDEND2), .Y(
        PARSETDEND2) );
    zan2b U399 ( .A(PER_CMDSTART1), .B(n1628), .Y(ICMDSTART1) );
    zan2b U400 ( .A(EHCI_MAC_EOT), .B(SITD_ACT1), .Y(SITD_MAC_EOT1) );
    zan2b U401 ( .A(EXESITD1), .B(n1680), .Y(SIPCIEND1) );
    zan2b U402 ( .A(PER_CMDSTART2), .B(n1631), .Y(QCMDSTART2) );
    zan2b U403 ( .A(n1680), .B(n1627), .Y(IPCIEND1) );
    zan2b U404 ( .A(EXESITD2), .B(n1679), .Y(SIPCIEND2) );
    zan2b U405 ( .A(EXESITD2), .B(PER_CMDSTART2), .Y(SICMDSTART2) );
    zao22b U406 ( .A(TDHCIGNT1), .B(n1681), .C(TDHCIGNT2), .D(n1682), .Y(
        HCIMWR) );
    zor3b U407 ( .A(IBUI_GO2), .B(QBUI_GO2), .C(SIBUI_GO2), .Y(BUI_GO2) );
    zan2b U408 ( .A(EXESITD2), .B(TD_PARSE_GO2), .Y(SITD_PARSE_GO2) );
    zan2b U409 ( .A(TD_PARSE_GO1), .B(n1637), .Y(ITD_PARSE_GO1) );
    zan2b U410 ( .A(EHCI_MAC_EOT), .B(ITD_ACT1), .Y(ITD_MAC_EOT1) );
    zor3b U411 ( .A(PARSESITDEND1), .B(PARSEITDEND1), .C(PARSEQHEND1), .Y(
        PARSETDEND1) );
    zan2b U412 ( .A(TD_PARSE_GO2), .B(n1639), .Y(ITD_PARSE_GO2) );
    zan2b U413 ( .A(n1680), .B(n1633), .Y(QPCIEND1) );
    zan2b U414 ( .A(EXESITD1), .B(TD_PARSE_GO1), .Y(SITD_PARSE_GO1) );
    zan2b U415 ( .A(EHCI_MAC_EOT), .B(ITD_ACT2), .Y(ITD_MAC_EOT2) );
    zor3b U416 ( .A(SICACHE_INVALID1), .B(ICACHE_INVALID1), .C(QCACHE_INVALID1
        ), .Y(CACHE_INVALID1) );
    zor3b U417 ( .A(IHCIREQ1), .B(QHCIREQ1), .C(SIHCIREQ1), .Y(TDHCIREQ1) );
    zor3b U418 ( .A(IEOT2), .B(QEOT2), .C(SIEOT2), .Y(EOT2) );
    zan2b U419 ( .A(n1679), .B(n1631), .Y(QPCIEND2) );
    zor3b U420 ( .A(ITDPARSING2), .B(QHPARSING2), .C(SITDPARSING2), .Y(
        TDPARSING2) );
    zan2b U421 ( .A(EXESITD1), .B(PER_CMDSTART1), .Y(SICMDSTART1) );
    zor3b U422 ( .A(ICMDSTART_REQ1), .B(QCMDSTART_REQ1), .C(SICMDSTART_REQ1), 
        .Y(PER_CMDSTART_REQ1) );
    zor3b U423 ( .A(IEOT1), .B(QEOT1), .C(SIEOT1), .Y(EOT1) );
    zan2b U424 ( .A(TD_ACT2), .B(EXESITD2), .Y(SITD_ACT2) );
    zan2b U425 ( .A(TD_ACT1), .B(EXESITD1), .Y(SITD_ACT1) );
    zan2b U426 ( .A(TDHCIGNT2), .B(PCIEND), .Y(n1679) );
    zan2b U427 ( .A(TDHCIGNT1), .B(PCIEND), .Y(n1680) );
    zan2b U428 ( .A(TD_ACT2), .B(n1631), .Y(QH_ACT2) );
    zan2b U429 ( .A(TD_ACT1), .B(n1633), .Y(QH_ACT1) );
    zan2b U430 ( .A(TD_ACT2), .B(n1626), .Y(ITD_ACT2) );
    zan2b U431 ( .A(TD_ACT1), .B(n1636), .Y(ITD_ACT1) );
    znr2b U432 ( .A(TD_CACHE_EN2), .B(TD_CACHE_EN1), .Y(n1669) );
    zinr2b U433 ( .A(TD_CACHE_EN2), .B(TD_CACHE_EN1), .Y(n1667) );
    znr2b U434 ( .A(TDHCIGNT2), .B(TDHCIGNT1), .Y(n1659) );
    zinr2b U435 ( .A(TDHCIGNT2), .B(TDHCIGNT1), .Y(n1657) );
    zmux21hb U436 ( .A(SIUP_LDW2_3), .B(QUP_LDW2_3), .S(n1632), .Y(UP_LDW2_3)
         );
    zmux21hb U437 ( .A(SIUP_LDW1_3), .B(QUP_LDW1_3), .S(n1634), .Y(UP_LDW1_3)
         );
    zmux21hb U438 ( .A(SIUP_DW2_3[9]), .B(QUP_DW2_3[9]), .S(n1631), .Y(
        UP_DW2_3[9]) );
    zmux21hb U439 ( .A(SIUP_DW2_3[8]), .B(QUP_DW2_3[8]), .S(n1632), .Y(
        UP_DW2_3[8]) );
    zmux21hb U440 ( .A(SIUP_DW2_3[7]), .B(QUP_DW2_3[7]), .S(n1631), .Y(
        UP_DW2_3[7]) );
    zmux21hb U441 ( .A(SIUP_DW2_3[6]), .B(QUP_DW2_3[6]), .S(n1632), .Y(
        UP_DW2_3[6]) );
    zmux21hb U442 ( .A(SIUP_DW2_3[5]), .B(QUP_DW2_3[5]), .S(n1631), .Y(
        UP_DW2_3[5]) );
    zmux21hb U443 ( .A(SIUP_DW2_3[4]), .B(QUP_DW2_3[4]), .S(n1632), .Y(
        UP_DW2_3[4]) );
    zmux21hb U444 ( .A(SIUP_DW2_3[31]), .B(QUP_DW2_3[31]), .S(n1631), .Y(
        UP_DW2_3[31]) );
    zmux21hb U445 ( .A(SIUP_DW2_3[30]), .B(QUP_DW2_3[30]), .S(n1632), .Y(
        UP_DW2_3[30]) );
    zmux21hb U446 ( .A(SIUP_DW2_3[3]), .B(QUP_DW2_3[3]), .S(n1631), .Y(
        UP_DW2_3[3]) );
    zmux21hb U447 ( .A(SIUP_DW2_3[29]), .B(QUP_DW2_3[29]), .S(n1632), .Y(
        UP_DW2_3[29]) );
    zmux21hb U448 ( .A(SIUP_DW2_3[28]), .B(QUP_DW2_3[28]), .S(n1631), .Y(
        UP_DW2_3[28]) );
    zmux21hb U449 ( .A(SIUP_DW2_3[27]), .B(QUP_DW2_3[27]), .S(n1632), .Y(
        UP_DW2_3[27]) );
    zmux21hb U450 ( .A(SIUP_DW2_3[26]), .B(QUP_DW2_3[26]), .S(n1631), .Y(
        UP_DW2_3[26]) );
    zmux21hb U451 ( .A(SIUP_DW2_3[25]), .B(QUP_DW2_3[25]), .S(n1632), .Y(
        UP_DW2_3[25]) );
    zmux21hb U452 ( .A(SIUP_DW2_3[24]), .B(QUP_DW2_3[24]), .S(n1632), .Y(
        UP_DW2_3[24]) );
    zmux21hb U453 ( .A(SIUP_DW2_3[23]), .B(QUP_DW2_3[23]), .S(n1632), .Y(
        UP_DW2_3[23]) );
    zmux21hb U454 ( .A(SIUP_DW2_3[22]), .B(QUP_DW2_3[22]), .S(n1632), .Y(
        UP_DW2_3[22]) );
    zmux21hb U455 ( .A(SIUP_DW2_3[21]), .B(QUP_DW2_3[21]), .S(n1632), .Y(
        UP_DW2_3[21]) );
    zmux21hb U456 ( .A(SIUP_DW2_3[20]), .B(QUP_DW2_3[20]), .S(n1632), .Y(
        UP_DW2_3[20]) );
    zmux21hb U457 ( .A(SIUP_DW2_3[2]), .B(QUP_DW2_3[2]), .S(n1632), .Y(
        UP_DW2_3[2]) );
    zmux21hb U458 ( .A(SIUP_DW2_3[19]), .B(QUP_DW2_3[19]), .S(n1632), .Y(
        UP_DW2_3[19]) );
    zmux21hb U459 ( .A(SIUP_DW2_3[18]), .B(QUP_DW2_3[18]), .S(n1632), .Y(
        UP_DW2_3[18]) );
    zmux21hb U460 ( .A(SIUP_DW2_3[17]), .B(QUP_DW2_3[17]), .S(n1632), .Y(
        UP_DW2_3[17]) );
    zmux21hb U461 ( .A(SIUP_DW2_3[16]), .B(QUP_DW2_3[16]), .S(n1632), .Y(
        UP_DW2_3[16]) );
    zmux21hb U462 ( .A(SIUP_DW2_3[15]), .B(QUP_DW2_3[15]), .S(n1632), .Y(
        UP_DW2_3[15]) );
    zmux21hb U463 ( .A(SIUP_DW2_3[14]), .B(QUP_DW2_3[14]), .S(n1631), .Y(
        UP_DW2_3[14]) );
    zmux21hb U464 ( .A(SIUP_DW2_3[13]), .B(QUP_DW2_3[13]), .S(n1631), .Y(
        UP_DW2_3[13]) );
    zmux21hb U465 ( .A(SIUP_DW2_3[12]), .B(QUP_DW2_3[12]), .S(n1631), .Y(
        UP_DW2_3[12]) );
    zmux21hb U466 ( .A(SIUP_DW2_3[11]), .B(QUP_DW2_3[11]), .S(n1631), .Y(
        UP_DW2_3[11]) );
    zmux21hb U467 ( .A(SIUP_DW2_3[10]), .B(QUP_DW2_3[10]), .S(n1631), .Y(
        UP_DW2_3[10]) );
    zmux21hb U468 ( .A(SIUP_DW2_3[1]), .B(QUP_DW2_3[1]), .S(n1631), .Y(
        UP_DW2_3[1]) );
    zmux21hb U469 ( .A(SIUP_DW2_3[0]), .B(QUP_DW2_3[0]), .S(n1631), .Y(
        UP_DW2_3[0]) );
    zmux21hb U470 ( .A(SIUP_DW1_3[9]), .B(QUP_DW1_3[9]), .S(n1633), .Y(
        UP_DW1_3[9]) );
    zmux21hb U471 ( .A(SIUP_DW1_3[8]), .B(QUP_DW1_3[8]), .S(n1634), .Y(
        UP_DW1_3[8]) );
    zmux21hb U472 ( .A(SIUP_DW1_3[7]), .B(QUP_DW1_3[7]), .S(n1633), .Y(
        UP_DW1_3[7]) );
    zmux21hb U473 ( .A(SIUP_DW1_3[6]), .B(QUP_DW1_3[6]), .S(n1634), .Y(
        UP_DW1_3[6]) );
    zmux21hb U474 ( .A(SIUP_DW1_3[5]), .B(QUP_DW1_3[5]), .S(n1633), .Y(
        UP_DW1_3[5]) );
    zmux21hb U475 ( .A(SIUP_DW1_3[4]), .B(QUP_DW1_3[4]), .S(n1634), .Y(
        UP_DW1_3[4]) );
    zmux21hb U476 ( .A(SIUP_DW1_3[31]), .B(QUP_DW1_3[31]), .S(n1633), .Y(
        UP_DW1_3[31]) );
    zmux21hb U477 ( .A(SIUP_DW1_3[30]), .B(QUP_DW1_3[30]), .S(n1634), .Y(
        UP_DW1_3[30]) );
    zmux21hb U478 ( .A(SIUP_DW1_3[3]), .B(QUP_DW1_3[3]), .S(n1633), .Y(
        UP_DW1_3[3]) );
    zmux21hb U479 ( .A(SIUP_DW1_3[29]), .B(QUP_DW1_3[29]), .S(n1634), .Y(
        UP_DW1_3[29]) );
    zmux21hb U480 ( .A(SIUP_DW1_3[28]), .B(QUP_DW1_3[28]), .S(n1633), .Y(
        UP_DW1_3[28]) );
    zmux21hb U481 ( .A(SIUP_DW1_3[27]), .B(QUP_DW1_3[27]), .S(n1634), .Y(
        UP_DW1_3[27]) );
    zmux21hb U482 ( .A(SIUP_DW1_3[26]), .B(QUP_DW1_3[26]), .S(n1633), .Y(
        UP_DW1_3[26]) );
    zmux21hb U483 ( .A(SIUP_DW1_3[25]), .B(QUP_DW1_3[25]), .S(n1634), .Y(
        UP_DW1_3[25]) );
    zmux21hb U484 ( .A(SIUP_DW1_3[24]), .B(QUP_DW1_3[24]), .S(n1634), .Y(
        UP_DW1_3[24]) );
    zmux21hb U485 ( .A(SIUP_DW1_3[23]), .B(QUP_DW1_3[23]), .S(n1634), .Y(
        UP_DW1_3[23]) );
    zmux21hb U486 ( .A(SIUP_DW1_3[22]), .B(QUP_DW1_3[22]), .S(n1634), .Y(
        UP_DW1_3[22]) );
    zmux21hb U487 ( .A(SIUP_DW1_3[21]), .B(QUP_DW1_3[21]), .S(n1634), .Y(
        UP_DW1_3[21]) );
    zmux21hb U488 ( .A(SIUP_DW1_3[20]), .B(QUP_DW1_3[20]), .S(n1634), .Y(
        UP_DW1_3[20]) );
    zmux21hb U489 ( .A(SIUP_DW1_3[2]), .B(QUP_DW1_3[2]), .S(n1634), .Y(
        UP_DW1_3[2]) );
    zmux21hb U490 ( .A(SIUP_DW1_3[19]), .B(QUP_DW1_3[19]), .S(n1634), .Y(
        UP_DW1_3[19]) );
    zmux21hb U491 ( .A(SIUP_DW1_3[18]), .B(QUP_DW1_3[18]), .S(n1634), .Y(
        UP_DW1_3[18]) );
    zmux21hb U492 ( .A(SIUP_DW1_3[17]), .B(QUP_DW1_3[17]), .S(n1634), .Y(
        UP_DW1_3[17]) );
    zmux21hb U493 ( .A(SIUP_DW1_3[16]), .B(QUP_DW1_3[16]), .S(n1634), .Y(
        UP_DW1_3[16]) );
    zmux21hb U494 ( .A(SIUP_DW1_3[15]), .B(QUP_DW1_3[15]), .S(n1634), .Y(
        UP_DW1_3[15]) );
    zmux21hb U495 ( .A(SIUP_DW1_3[14]), .B(QUP_DW1_3[14]), .S(n1633), .Y(
        UP_DW1_3[14]) );
    zmux21hb U496 ( .A(SIUP_DW1_3[13]), .B(QUP_DW1_3[13]), .S(n1633), .Y(
        UP_DW1_3[13]) );
    zmux21hb U497 ( .A(SIUP_DW1_3[12]), .B(QUP_DW1_3[12]), .S(n1633), .Y(
        UP_DW1_3[12]) );
    zmux21hb U498 ( .A(SIUP_DW1_3[11]), .B(QUP_DW1_3[11]), .S(n1633), .Y(
        UP_DW1_3[11]) );
    zmux21hb U499 ( .A(SIUP_DW1_3[10]), .B(QUP_DW1_3[10]), .S(n1633), .Y(
        UP_DW1_3[10]) );
    zmux21hb U500 ( .A(SIUP_DW1_3[1]), .B(QUP_DW1_3[1]), .S(n1633), .Y(
        UP_DW1_3[1]) );
    zmux21hb U501 ( .A(SIUP_DW1_3[0]), .B(QUP_DW1_3[0]), .S(n1633), .Y(
        UP_DW1_3[0]) );
    zmux21hb U502 ( .A(SICACHEPHASE2), .B(QCACHEPHASE2), .S(n1631), .Y(
        CACHEPHASE2) );
    zmux21hb U503 ( .A(SICACHEPHASE1), .B(QCACHEPHASE1), .S(n1633), .Y(
        CACHEPHASE1) );
    zao222b U504 ( .A(IMWR1), .B(n1637), .C(SIMWR1), .D(EXESITD1), .E(QHMWR1), 
        .F(n1633), .Y(n1681) );
    zao222b U505 ( .A(IMWR2), .B(n1639), .C(SIMWR2), .D(EXESITD2), .E(QHMWR2), 
        .F(n1631), .Y(n1682) );
    zao222b U506 ( .A(SIDWOFFSET2[3]), .B(n1646), .C(QHDWOFFSET2[3]), .D(n1653
        ), .E(IDWOFFSET2[3]), .F(n1640), .Y(n1675) );
    zao222b U507 ( .A(SIDWOFFSET1[3]), .B(n1643), .C(QHDWOFFSET1[3]), .D(n1648
        ), .E(IDWOFFSET1[3]), .F(n1627), .Y(n1676) );
    zao222b U508 ( .A(SIDWOFFSET2[2]), .B(n1619), .C(QHDWOFFSET2[2]), .D(n1654
        ), .E(IDWOFFSET2[2]), .F(n1626), .Y(n1673) );
    zao222b U509 ( .A(SIDWOFFSET1[2]), .B(n1623), .C(QHDWOFFSET1[2]), .D(n1649
        ), .E(IDWOFFSET1[2]), .F(n1628), .Y(n1674) );
    zao222b U510 ( .A(SIDWOFFSET2[1]), .B(n1610), .C(QHDWOFFSET2[1]), .D(n1622
        ), .E(IDWOFFSET2[1]), .F(n1626), .Y(n1671) );
    zao222b U511 ( .A(SIDWOFFSET1[1]), .B(n1612), .C(QHDWOFFSET1[1]), .D(n1618
        ), .E(IDWOFFSET1[1]), .F(n1636), .Y(n1672) );
    zao222b U512 ( .A(SIDWOFFSET2[0]), .B(n1645), .C(QHDWOFFSET2[0]), .D(n1653
        ), .E(IDWOFFSET2[0]), .F(n1640), .Y(n1668) );
    zao222b U513 ( .A(SIDWOFFSET1[0]), .B(n1642), .C(QHDWOFFSET1[0]), .D(n1648
        ), .E(IDWOFFSET1[0]), .F(n1627), .Y(n1670) );
    zao222b U514 ( .A(SIDWNUM2[3]), .B(n1644), .C(QHDWNUM2[3]), .D(n1654), .E(
        IDWNUM2[3]), .F(n1639), .Y(n1665) );
    zao222b U515 ( .A(SIDWNUM1[3]), .B(n1641), .C(QHDWNUM1[3]), .D(n1649), .E(
        IDWNUM1[3]), .F(n1635), .Y(n1666) );
    zao222b U516 ( .A(SIDWNUM2[2]), .B(n1646), .C(QHDWNUM2[2]), .D(n1653), .E(
        IDWNUM2[2]), .F(n1638), .Y(n1663) );
    zao222b U517 ( .A(SIDWNUM1[2]), .B(n1643), .C(QHDWNUM1[2]), .D(n1648), .E(
        IDWNUM1[2]), .F(n1637), .Y(n1664) );
    zao222b U518 ( .A(SIDWNUM2[1]), .B(n1610), .C(QHDWNUM2[1]), .D(n1655), .E(
        IDWNUM2[1]), .F(n1639), .Y(n1661) );
    zao222b U519 ( .A(SIDWNUM1[1]), .B(n1612), .C(QHDWNUM1[1]), .D(n1650), .E(
        IDWNUM1[1]), .F(n1635), .Y(n1662) );
    zao222b U520 ( .A(SIDWNUM2[0]), .B(n1644), .C(QHDWNUM2[0]), .D(n1622), .E(
        IDWNUM2[0]), .F(n1626), .Y(n1658) );
    zao222b U521 ( .A(SIDWNUM1[0]), .B(n1641), .C(QHDWNUM1[0]), .D(n1618), .E(
        IDWNUM1[0]), .F(n1636), .Y(n1660) );
endmodule


module PERIODIC_ADCTL ( PCICLK, TRST_, DWCNT, RUN, ADI, PERHCIADR, TDHCIGNT1, 
    TDHCIGNT2, EXEITD1, EXEITD2, EXESITD1, EXESITD2, IHCIADR1, IHCIADR2, 
    QHCIADR1, QHCIADR2, SIHCIADR1, SIHCIADR2, HCIADR, IHCIADD1, IHCIADD2, 
    QHCIADD1, QHCIADD2, SIHCIADD1, SIHCIADD2, HCIADD );
input  [3:0] DWCNT;
input  [31:0] ADI;
input  [31:0] IHCIADD2;
input  [31:0] QHCIADD1;
input  [31:0] SIHCIADD2;
input  [31:0] IHCIADR2;
input  [31:0] QHCIADR1;
input  [31:0] SIHCIADR2;
input  [31:0] PERHCIADR;
input  [31:0] IHCIADR1;
output [31:0] HCIADR;
input  [31:0] QHCIADD2;
input  [31:0] SIHCIADD1;
output [31:0] HCIADD;
input  [31:0] IHCIADD1;
input  [31:0] QHCIADR2;
input  [31:0] SIHCIADR1;
input  PCICLK, TRST_, RUN, TDHCIGNT1, TDHCIGNT2, EXEITD1, EXEITD2, EXESITD1, 
    EXESITD2;
    wire HCIADR_p_2, HCIADR_p_13, HCIADR_p_26, HCIADR_p_21, HCIADR_p_14, 
        HCIADR_p_5, HCIADR_p_28, HCIADR_p_20, HCIADR_p_29, HCIADR_p_4, 
        HCIADR_p_15, HCIADR_p_12, HCIADR_p_3, HCIADR_p_27, HCIADR_p_1, 
        HCIADR_p_10, HCIADR_p_25, HCIADR_p_8, HCIADR_p_19, HCIADR_p_22, 
        HCIADR_p_17, HCIADR_p_6, HCIADR_p_23, HCIADR_p_7, HCIADR_p_16, 
        HCIADR_p_11, HCIADR_p_0, HCIADR_p_18, HCIADR_p_9, HCIADR_p_24, 
        add_52_carry_29, add_52_carry_1, add_52_carry_20, add_52_carry_15, 
        add_52_carry_8, add_52_carry_28, add_52_carry_27, add_52_carry_26, 
        add_52_carry_12, add_52_carry_6, add_52_carry_14, add_52_carry_13, 
        add_52_carry_7, add_52_carry_24, add_52_carry_23, add_52_carry_21, 
        add_52_carry_16, add_52_carry_9, add_52_carry_2, add_52_carry_18, 
        add_52_carry_25, add_52_carry_11, add_52_carry_5, add_52_carry_19, 
        add_52_carry_10, add_52_carry_4, add_52_carry_22, add_52_carry_17, 
        add_52_carry_3, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
        n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, 
        n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
        n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
        n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, 
        n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, 
        n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, 
        n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, 
        n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, 
        n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
        n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
        n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
        n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
        n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
        n326, n327, n328, n329, n330, n331, n332, n333;
    assign HCIADR[1] = 1'b0;
    assign HCIADR[0] = 1'b0;
    zor2b U13 ( .A(n285), .B(n291), .Y(n307) );
    zor2b U14 ( .A(n285), .B(n286), .Y(n305) );
    zor2b U15 ( .A(EXEITD2), .B(EXESITD2), .Y(n286) );
    zor2b U16 ( .A(n285), .B(n289), .Y(n306) );
    zor2b U17 ( .A(EXEITD2), .B(n288), .Y(n289) );
    zivb U18 ( .A(EXESITD2), .Y(n288) );
    zor2b U19 ( .A(n293), .B(n299), .Y(n304) );
    zor2b U20 ( .A(n293), .B(n294), .Y(n302) );
    zor2b U21 ( .A(EXEITD1), .B(EXESITD1), .Y(n294) );
    zor2b U22 ( .A(n293), .B(n297), .Y(n303) );
    zor2b U23 ( .A(EXEITD1), .B(n296), .Y(n297) );
    zivb U24 ( .A(EXESITD1), .Y(n296) );
    zaoi2x4b U25 ( .A(QHCIADR2[2]), .B(n308), .C(SIHCIADR2[2]), .D(n309), .E(
        IHCIADR2[2]), .F(n310), .G(QHCIADR1[2]), .H(n311), .Y(n226) );
    zaoi2x4b U26 ( .A(QHCIADR2[3]), .B(n330), .C(SIHCIADR2[3]), .D(n331), .E(
        IHCIADR2[3]), .F(n332), .G(QHCIADR1[3]), .H(n333), .Y(n228) );
    zaoi2x4b U27 ( .A(QHCIADR2[4]), .B(n308), .C(SIHCIADR2[4]), .D(n309), .E(
        IHCIADR2[4]), .F(n310), .G(QHCIADR1[4]), .H(n311), .Y(n230) );
    zaoi2x4b U28 ( .A(QHCIADR2[5]), .B(n330), .C(SIHCIADR2[5]), .D(n331), .E(
        IHCIADR2[5]), .F(n332), .G(QHCIADR1[5]), .H(n333), .Y(n232) );
    zaoi2x4b U29 ( .A(QHCIADR2[6]), .B(n308), .C(SIHCIADR2[6]), .D(n309), .E(
        IHCIADR2[6]), .F(n310), .G(QHCIADR1[6]), .H(n311), .Y(n234) );
    zaoi2x4b U30 ( .A(QHCIADR2[7]), .B(n330), .C(SIHCIADR2[7]), .D(n331), .E(
        IHCIADR2[7]), .F(n332), .G(QHCIADR1[7]), .H(n333), .Y(n236) );
    zaoi2x4b U31 ( .A(QHCIADR2[8]), .B(n308), .C(SIHCIADR2[8]), .D(n309), .E(
        IHCIADR2[8]), .F(n310), .G(QHCIADR1[8]), .H(n311), .Y(n238) );
    zaoi2x4b U32 ( .A(QHCIADR2[9]), .B(n330), .C(SIHCIADR2[9]), .D(n331), .E(
        IHCIADR2[9]), .F(n332), .G(QHCIADR1[9]), .H(n333), .Y(n240) );
    zaoi2x4b U33 ( .A(QHCIADR2[10]), .B(n308), .C(SIHCIADR2[10]), .D(n309), 
        .E(IHCIADR2[10]), .F(n310), .G(QHCIADR1[10]), .H(n311), .Y(n242) );
    zaoi2x4b U34 ( .A(QHCIADR2[11]), .B(n330), .C(SIHCIADR2[11]), .D(n331), 
        .E(IHCIADR2[11]), .F(n332), .G(QHCIADR1[11]), .H(n333), .Y(n244) );
    zaoi2x4b U35 ( .A(QHCIADR2[12]), .B(n308), .C(SIHCIADR2[12]), .D(n309), 
        .E(IHCIADR2[12]), .F(n310), .G(QHCIADR1[12]), .H(n311), .Y(n246) );
    zaoi2x4b U36 ( .A(QHCIADR2[13]), .B(n330), .C(SIHCIADR2[13]), .D(n331), 
        .E(IHCIADR2[13]), .F(n332), .G(QHCIADR1[13]), .H(n333), .Y(n248) );
    zaoi2x4b U37 ( .A(QHCIADR2[14]), .B(n308), .C(SIHCIADR2[14]), .D(n309), 
        .E(IHCIADR2[14]), .F(n310), .G(QHCIADR1[14]), .H(n311), .Y(n250) );
    zaoi2x4b U38 ( .A(QHCIADR2[15]), .B(n330), .C(SIHCIADR2[15]), .D(n331), 
        .E(IHCIADR2[15]), .F(n332), .G(QHCIADR1[15]), .H(n333), .Y(n252) );
    zaoi2x4b U39 ( .A(QHCIADR2[16]), .B(n308), .C(SIHCIADR2[16]), .D(n309), 
        .E(IHCIADR2[16]), .F(n310), .G(QHCIADR1[16]), .H(n311), .Y(n254) );
    zaoi2x4b U40 ( .A(QHCIADR2[17]), .B(n330), .C(SIHCIADR2[17]), .D(n331), 
        .E(IHCIADR2[17]), .F(n332), .G(QHCIADR1[17]), .H(n333), .Y(n256) );
    zaoi2x4b U41 ( .A(QHCIADR2[18]), .B(n308), .C(SIHCIADR2[18]), .D(n309), 
        .E(IHCIADR2[18]), .F(n310), .G(QHCIADR1[18]), .H(n311), .Y(n258) );
    zaoi2x4b U42 ( .A(QHCIADR2[19]), .B(n330), .C(SIHCIADR2[19]), .D(n331), 
        .E(IHCIADR2[19]), .F(n332), .G(QHCIADR1[19]), .H(n333), .Y(n260) );
    zaoi2x4b U43 ( .A(QHCIADR2[20]), .B(n308), .C(SIHCIADR2[20]), .D(n309), 
        .E(IHCIADR2[20]), .F(n310), .G(QHCIADR1[20]), .H(n311), .Y(n262) );
    zaoi2x4b U44 ( .A(QHCIADR2[21]), .B(n330), .C(SIHCIADR2[21]), .D(n331), 
        .E(IHCIADR2[21]), .F(n332), .G(QHCIADR1[21]), .H(n333), .Y(n264) );
    zaoi2x4b U45 ( .A(QHCIADR2[22]), .B(n330), .C(SIHCIADR2[22]), .D(n331), 
        .E(IHCIADR2[22]), .F(n332), .G(QHCIADR1[22]), .H(n333), .Y(n266) );
    zaoi2x4b U46 ( .A(QHCIADR2[23]), .B(n308), .C(SIHCIADR2[23]), .D(n309), 
        .E(IHCIADR2[23]), .F(n310), .G(QHCIADR1[23]), .H(n311), .Y(n268) );
    zaoi2x4b U47 ( .A(QHCIADR2[24]), .B(n330), .C(SIHCIADR2[24]), .D(n331), 
        .E(IHCIADR2[24]), .F(n332), .G(QHCIADR1[24]), .H(n333), .Y(n270) );
    zaoi2x4b U48 ( .A(QHCIADR2[25]), .B(n308), .C(SIHCIADR2[25]), .D(n309), 
        .E(IHCIADR2[25]), .F(n310), .G(QHCIADR1[25]), .H(n311), .Y(n272) );
    zaoi2x4b U49 ( .A(QHCIADR2[26]), .B(n330), .C(SIHCIADR2[26]), .D(n331), 
        .E(IHCIADR2[26]), .F(n332), .G(QHCIADR1[26]), .H(n333), .Y(n274) );
    zaoi2x4b U50 ( .A(QHCIADR2[27]), .B(n308), .C(SIHCIADR2[27]), .D(n309), 
        .E(IHCIADR2[27]), .F(n310), .G(QHCIADR1[27]), .H(n311), .Y(n276) );
    zaoi2x4b U51 ( .A(QHCIADR2[28]), .B(n330), .C(SIHCIADR2[28]), .D(n331), 
        .E(IHCIADR2[28]), .F(n332), .G(QHCIADR1[28]), .H(n333), .Y(n278) );
    zaoi2x4b U52 ( .A(QHCIADR2[29]), .B(n308), .C(SIHCIADR2[29]), .D(n309), 
        .E(IHCIADR2[29]), .F(n310), .G(QHCIADR1[29]), .H(n311), .Y(n280) );
    zaoi2x4b U53 ( .A(QHCIADR2[30]), .B(n330), .C(SIHCIADR2[30]), .D(n331), 
        .E(IHCIADR2[30]), .F(n332), .G(QHCIADR1[30]), .H(n333), .Y(n282) );
    zaoi2x4b U54 ( .A(QHCIADR2[31]), .B(n308), .C(SIHCIADR2[31]), .D(n309), 
        .E(IHCIADR2[31]), .F(n310), .G(QHCIADR1[31]), .H(n311), .Y(n284) );
    zivc U55 ( .A(n287), .Y(n308) );
    zor2b U56 ( .A(n285), .B(n286), .Y(n287) );
    zivb U57 ( .A(TDHCIGNT2), .Y(n285) );
    zivc U58 ( .A(n290), .Y(n309) );
    zor2b U59 ( .A(n285), .B(n289), .Y(n290) );
    zivc U60 ( .A(n292), .Y(n310) );
    zor2b U61 ( .A(n285), .B(n291), .Y(n292) );
    zivb U62 ( .A(EXEITD2), .Y(n291) );
    zivc U63 ( .A(n295), .Y(n311) );
    zor2b U64 ( .A(n293), .B(n294), .Y(n295) );
    zivc U65 ( .A(n287), .Y(n330) );
    zivc U66 ( .A(n290), .Y(n331) );
    zivc U67 ( .A(n292), .Y(n332) );
    zivc U68 ( .A(n295), .Y(n333) );
    zivc U69 ( .A(n300), .Y(n312) );
    zor2b U70 ( .A(n293), .B(n299), .Y(n300) );
    zivb U71 ( .A(TDHCIGNT1), .Y(n293) );
    zivb U72 ( .A(EXEITD1), .Y(n299) );
    zivc U73 ( .A(n301), .Y(n328) );
    zor2b U74 ( .A(TDHCIGNT2), .B(TDHCIGNT1), .Y(n301) );
    zivc U75 ( .A(n298), .Y(n314) );
    zor2b U76 ( .A(n293), .B(n297), .Y(n298) );
    zivc U77 ( .A(n300), .Y(n327) );
    zivc U78 ( .A(n301), .Y(n313) );
    zivc U79 ( .A(n298), .Y(n329) );
    zor2b U80 ( .A(n219), .B(n220), .Y(HCIADD[0]) );
    zor2b U81 ( .A(n215), .B(n216), .Y(HCIADD[1]) );
    zor2b U82 ( .A(n201), .B(n202), .Y(HCIADD[2]) );
    zor2b U83 ( .A(n173), .B(n174), .Y(HCIADD[3]) );
    zor2b U84 ( .A(n183), .B(n184), .Y(HCIADD[4]) );
    zor2b U85 ( .A(n203), .B(n204), .Y(HCIADD[5]) );
    zor2b U86 ( .A(n211), .B(n212), .Y(HCIADD[6]) );
    zor2b U87 ( .A(n195), .B(n196), .Y(HCIADD[7]) );
    zor2b U88 ( .A(n223), .B(n224), .Y(HCIADD[8]) );
    zor2b U89 ( .A(n189), .B(n190), .Y(HCIADD[9]) );
    zor2b U90 ( .A(n165), .B(n166), .Y(HCIADD[10]) );
    zor2b U91 ( .A(n171), .B(n172), .Y(HCIADD[11]) );
    zor2b U92 ( .A(n177), .B(n178), .Y(HCIADD[12]) );
    zor2b U93 ( .A(n207), .B(n208), .Y(HCIADD[13]) );
    zor2b U94 ( .A(n199), .B(n200), .Y(HCIADD[14]) );
    zor2b U95 ( .A(n187), .B(n188), .Y(HCIADD[15]) );
    zor2b U96 ( .A(n163), .B(n164), .Y(HCIADD[16]) );
    zor2b U97 ( .A(n181), .B(n182), .Y(HCIADD[17]) );
    zor2b U98 ( .A(n175), .B(n176), .Y(HCIADD[18]) );
    zor2b U99 ( .A(n205), .B(n206), .Y(HCIADD[19]) );
    zor2b U100 ( .A(n213), .B(n214), .Y(HCIADD[20]) );
    zor2b U101 ( .A(n221), .B(n222), .Y(HCIADD[21]) );
    zor2b U102 ( .A(n191), .B(n192), .Y(HCIADD[22]) );
    zor2b U103 ( .A(n161), .B(n162), .Y(HCIADD[23]) );
    zor2b U104 ( .A(n185), .B(n186), .Y(HCIADD[24]) );
    zor2b U105 ( .A(n193), .B(n194), .Y(HCIADD[25]) );
    zor2b U106 ( .A(n217), .B(n218), .Y(HCIADD[26]) );
    zor2b U107 ( .A(n197), .B(n198), .Y(HCIADD[27]) );
    zor2b U108 ( .A(n209), .B(n210), .Y(HCIADD[28]) );
    zor2b U109 ( .A(n179), .B(n180), .Y(HCIADD[29]) );
    zor2b U110 ( .A(n169), .B(n170), .Y(HCIADD[30]) );
    zivc U111 ( .A(n303), .Y(n315) );
    zivc U112 ( .A(n302), .Y(n316) );
    zivc U113 ( .A(n304), .Y(n317) );
    zivc U114 ( .A(n306), .Y(n318) );
    zivc U115 ( .A(n305), .Y(n319) );
    zivc U116 ( .A(n307), .Y(n320) );
    zor2b U117 ( .A(n167), .B(n168), .Y(HCIADD[31]) );
    zivc U118 ( .A(n303), .Y(n321) );
    zivc U119 ( .A(n302), .Y(n322) );
    zivc U120 ( .A(n304), .Y(n323) );
    zivc U121 ( .A(n306), .Y(n324) );
    zivc U122 ( .A(n305), .Y(n325) );
    zivc U123 ( .A(n307), .Y(n326) );
    zxo2b U124 ( .A(add_52_carry_29), .B(HCIADR_p_29), .Y(HCIADR[31]) );
    zan2b U125 ( .A(HCIADR_p_28), .B(add_52_carry_28), .Y(add_52_carry_29) );
    zxo2b U126 ( .A(HCIADR_p_28), .B(add_52_carry_28), .Y(HCIADR[30]) );
    zan2b U127 ( .A(HCIADR_p_27), .B(add_52_carry_27), .Y(add_52_carry_28) );
    zxo2b U128 ( .A(HCIADR_p_27), .B(add_52_carry_27), .Y(HCIADR[29]) );
    zan2b U129 ( .A(HCIADR_p_26), .B(add_52_carry_26), .Y(add_52_carry_27) );
    zxo2b U130 ( .A(HCIADR_p_26), .B(add_52_carry_26), .Y(HCIADR[28]) );
    zan2b U131 ( .A(HCIADR_p_25), .B(add_52_carry_25), .Y(add_52_carry_26) );
    zxo2b U132 ( .A(HCIADR_p_25), .B(add_52_carry_25), .Y(HCIADR[27]) );
    zan2b U133 ( .A(HCIADR_p_24), .B(add_52_carry_24), .Y(add_52_carry_25) );
    zxo2b U134 ( .A(HCIADR_p_24), .B(add_52_carry_24), .Y(HCIADR[26]) );
    zan2b U135 ( .A(HCIADR_p_23), .B(add_52_carry_23), .Y(add_52_carry_24) );
    zxo2b U136 ( .A(HCIADR_p_23), .B(add_52_carry_23), .Y(HCIADR[25]) );
    zan2b U137 ( .A(HCIADR_p_22), .B(add_52_carry_22), .Y(add_52_carry_23) );
    zxo2b U138 ( .A(HCIADR_p_22), .B(add_52_carry_22), .Y(HCIADR[24]) );
    zan2b U139 ( .A(HCIADR_p_21), .B(add_52_carry_21), .Y(add_52_carry_22) );
    zxo2b U140 ( .A(HCIADR_p_21), .B(add_52_carry_21), .Y(HCIADR[23]) );
    zan2b U141 ( .A(HCIADR_p_20), .B(add_52_carry_20), .Y(add_52_carry_21) );
    zxo2b U142 ( .A(HCIADR_p_20), .B(add_52_carry_20), .Y(HCIADR[22]) );
    zan2b U143 ( .A(HCIADR_p_19), .B(add_52_carry_19), .Y(add_52_carry_20) );
    zxo2b U144 ( .A(HCIADR_p_19), .B(add_52_carry_19), .Y(HCIADR[21]) );
    zan2b U145 ( .A(HCIADR_p_18), .B(add_52_carry_18), .Y(add_52_carry_19) );
    zxo2b U146 ( .A(HCIADR_p_18), .B(add_52_carry_18), .Y(HCIADR[20]) );
    zan2b U147 ( .A(HCIADR_p_17), .B(add_52_carry_17), .Y(add_52_carry_18) );
    zxo2b U148 ( .A(HCIADR_p_17), .B(add_52_carry_17), .Y(HCIADR[19]) );
    zan2b U149 ( .A(HCIADR_p_16), .B(add_52_carry_16), .Y(add_52_carry_17) );
    zxo2b U150 ( .A(HCIADR_p_16), .B(add_52_carry_16), .Y(HCIADR[18]) );
    zan2b U151 ( .A(HCIADR_p_15), .B(add_52_carry_15), .Y(add_52_carry_16) );
    zxo2b U152 ( .A(HCIADR_p_15), .B(add_52_carry_15), .Y(HCIADR[17]) );
    zan2b U153 ( .A(HCIADR_p_14), .B(add_52_carry_14), .Y(add_52_carry_15) );
    zxo2b U154 ( .A(HCIADR_p_14), .B(add_52_carry_14), .Y(HCIADR[16]) );
    zan2b U155 ( .A(HCIADR_p_13), .B(add_52_carry_13), .Y(add_52_carry_14) );
    zxo2b U156 ( .A(HCIADR_p_13), .B(add_52_carry_13), .Y(HCIADR[15]) );
    zan2b U157 ( .A(HCIADR_p_12), .B(add_52_carry_12), .Y(add_52_carry_13) );
    zxo2b U158 ( .A(HCIADR_p_12), .B(add_52_carry_12), .Y(HCIADR[14]) );
    zan2b U159 ( .A(HCIADR_p_11), .B(add_52_carry_11), .Y(add_52_carry_12) );
    zxo2b U160 ( .A(HCIADR_p_11), .B(add_52_carry_11), .Y(HCIADR[13]) );
    zan2b U161 ( .A(HCIADR_p_10), .B(add_52_carry_10), .Y(add_52_carry_11) );
    zxo2b U162 ( .A(HCIADR_p_10), .B(add_52_carry_10), .Y(HCIADR[12]) );
    zan2b U163 ( .A(HCIADR_p_9), .B(add_52_carry_9), .Y(add_52_carry_10) );
    zxo2b U164 ( .A(HCIADR_p_9), .B(add_52_carry_9), .Y(HCIADR[11]) );
    zan2b U165 ( .A(HCIADR_p_8), .B(add_52_carry_8), .Y(add_52_carry_9) );
    zxo2b U166 ( .A(HCIADR_p_8), .B(add_52_carry_8), .Y(HCIADR[10]) );
    zan2b U167 ( .A(HCIADR_p_7), .B(add_52_carry_7), .Y(add_52_carry_8) );
    zxo2b U168 ( .A(HCIADR_p_7), .B(add_52_carry_7), .Y(HCIADR[9]) );
    zan2b U169 ( .A(HCIADR_p_6), .B(add_52_carry_6), .Y(add_52_carry_7) );
    zxo2b U170 ( .A(HCIADR_p_6), .B(add_52_carry_6), .Y(HCIADR[8]) );
    zan2b U171 ( .A(HCIADR_p_5), .B(add_52_carry_5), .Y(add_52_carry_6) );
    zxo2b U172 ( .A(HCIADR_p_5), .B(add_52_carry_5), .Y(HCIADR[7]) );
    zan2b U173 ( .A(HCIADR_p_4), .B(add_52_carry_4), .Y(add_52_carry_5) );
    zxo2b U174 ( .A(HCIADR_p_4), .B(add_52_carry_4), .Y(HCIADR[6]) );
    zan2b U175 ( .A(DWCNT[0]), .B(HCIADR_p_0), .Y(add_52_carry_1) );
    zxo2b U176 ( .A(DWCNT[0]), .B(HCIADR_p_0), .Y(HCIADR[2]) );
    zfa1b add_52_U1_3 ( .A(HCIADR_p_3), .B(DWCNT[3]), .CI(add_52_carry_3), 
        .CO(add_52_carry_4), .S(HCIADR[5]) );
    zfa1b add_52_U1_2 ( .A(HCIADR_p_2), .B(DWCNT[2]), .CI(add_52_carry_2), 
        .CO(add_52_carry_3), .S(HCIADR[4]) );
    zfa1b add_52_U1_1 ( .A(HCIADR_p_1), .B(DWCNT[1]), .CI(add_52_carry_1), 
        .CO(add_52_carry_2), .S(HCIADR[3]) );
    zind2d U177 ( .A(n225), .B(n226), .Y(HCIADR_p_0) );
    zind2d U178 ( .A(n227), .B(n228), .Y(HCIADR_p_1) );
    zind2d U179 ( .A(n229), .B(n230), .Y(HCIADR_p_2) );
    zind2d U180 ( .A(n231), .B(n232), .Y(HCIADR_p_3) );
    zind2d U181 ( .A(n233), .B(n234), .Y(HCIADR_p_4) );
    zind2d U182 ( .A(n235), .B(n236), .Y(HCIADR_p_5) );
    zind2d U183 ( .A(n237), .B(n238), .Y(HCIADR_p_6) );
    zind2d U184 ( .A(n239), .B(n240), .Y(HCIADR_p_7) );
    zind2d U185 ( .A(n241), .B(n242), .Y(HCIADR_p_8) );
    zind2d U186 ( .A(n243), .B(n244), .Y(HCIADR_p_9) );
    zind2d U187 ( .A(n245), .B(n246), .Y(HCIADR_p_10) );
    zind2d U188 ( .A(n247), .B(n248), .Y(HCIADR_p_11) );
    zind2d U189 ( .A(n249), .B(n250), .Y(HCIADR_p_12) );
    zind2d U190 ( .A(n251), .B(n252), .Y(HCIADR_p_13) );
    zind2d U191 ( .A(n253), .B(n254), .Y(HCIADR_p_14) );
    zind2d U192 ( .A(n255), .B(n256), .Y(HCIADR_p_15) );
    zind2d U193 ( .A(n257), .B(n258), .Y(HCIADR_p_16) );
    zind2d U194 ( .A(n259), .B(n260), .Y(HCIADR_p_17) );
    zind2d U195 ( .A(n261), .B(n262), .Y(HCIADR_p_18) );
    zind2d U196 ( .A(n263), .B(n264), .Y(HCIADR_p_19) );
    zind2d U197 ( .A(n265), .B(n266), .Y(HCIADR_p_20) );
    zind2d U198 ( .A(n267), .B(n268), .Y(HCIADR_p_21) );
    zind2d U199 ( .A(n269), .B(n270), .Y(HCIADR_p_22) );
    zind2d U200 ( .A(n271), .B(n272), .Y(HCIADR_p_23) );
    zind2d U201 ( .A(n273), .B(n274), .Y(HCIADR_p_24) );
    zind2d U202 ( .A(n275), .B(n276), .Y(HCIADR_p_25) );
    zind2d U203 ( .A(n277), .B(n278), .Y(HCIADR_p_26) );
    zind2d U204 ( .A(n279), .B(n280), .Y(HCIADR_p_27) );
    zind2d U205 ( .A(n281), .B(n282), .Y(HCIADR_p_28) );
    zind2d U206 ( .A(n283), .B(n284), .Y(HCIADR_p_29) );
    zao222b U207 ( .A(IHCIADR1[11]), .B(n327), .C(n313), .D(PERHCIADR[11]), 
        .E(SIHCIADR1[11]), .F(n329), .Y(n243) );
    zao222b U208 ( .A(IHCIADR1[10]), .B(n312), .C(PERHCIADR[10]), .D(n328), 
        .E(SIHCIADR1[10]), .F(n314), .Y(n241) );
    zao222b U209 ( .A(IHCIADR1[9]), .B(n327), .C(PERHCIADR[9]), .D(n313), .E(
        SIHCIADR1[9]), .F(n329), .Y(n239) );
    zao222b U210 ( .A(IHCIADR1[8]), .B(n312), .C(PERHCIADR[8]), .D(n328), .E(
        SIHCIADR1[8]), .F(n314), .Y(n237) );
    zao222b U211 ( .A(IHCIADR1[7]), .B(n327), .C(PERHCIADR[7]), .D(n313), .E(
        SIHCIADR1[7]), .F(n329), .Y(n235) );
    zao222b U212 ( .A(IHCIADR1[6]), .B(n312), .C(PERHCIADR[6]), .D(n328), .E(
        SIHCIADR1[6]), .F(n314), .Y(n233) );
    zao222b U213 ( .A(IHCIADR1[5]), .B(n327), .C(PERHCIADR[5]), .D(n313), .E(
        SIHCIADR1[5]), .F(n329), .Y(n231) );
    zao222b U214 ( .A(IHCIADR1[31]), .B(n312), .C(PERHCIADR[31]), .D(n328), 
        .E(SIHCIADR1[31]), .F(n314), .Y(n283) );
    zao222b U215 ( .A(IHCIADR1[30]), .B(n327), .C(PERHCIADR[30]), .D(n313), 
        .E(SIHCIADR1[30]), .F(n329), .Y(n281) );
    zao222b U216 ( .A(IHCIADR1[29]), .B(n312), .C(PERHCIADR[29]), .D(n328), 
        .E(SIHCIADR1[29]), .F(n314), .Y(n279) );
    zao222b U217 ( .A(IHCIADR1[28]), .B(n327), .C(PERHCIADR[28]), .D(n313), 
        .E(SIHCIADR1[28]), .F(n329), .Y(n277) );
    zao222b U218 ( .A(IHCIADR1[27]), .B(n312), .C(PERHCIADR[27]), .D(n328), 
        .E(SIHCIADR1[27]), .F(n314), .Y(n275) );
    zao222b U219 ( .A(IHCIADR1[26]), .B(n327), .C(PERHCIADR[26]), .D(n313), 
        .E(SIHCIADR1[26]), .F(n329), .Y(n273) );
    zao222b U220 ( .A(IHCIADR1[25]), .B(n312), .C(PERHCIADR[25]), .D(n328), 
        .E(SIHCIADR1[25]), .F(n314), .Y(n271) );
    zao222b U221 ( .A(IHCIADR1[24]), .B(n327), .C(PERHCIADR[24]), .D(n313), 
        .E(SIHCIADR1[24]), .F(n329), .Y(n269) );
    zao222b U222 ( .A(IHCIADR1[23]), .B(n312), .C(PERHCIADR[23]), .D(n328), 
        .E(SIHCIADR1[23]), .F(n314), .Y(n267) );
    zao222b U223 ( .A(IHCIADR1[22]), .B(n327), .C(PERHCIADR[22]), .D(n313), 
        .E(SIHCIADR1[22]), .F(n329), .Y(n265) );
    zao222b U224 ( .A(IHCIADR1[4]), .B(n312), .C(PERHCIADR[4]), .D(n328), .E(
        SIHCIADR1[4]), .F(n314), .Y(n229) );
    zao222b U225 ( .A(IHCIADR1[21]), .B(n327), .C(PERHCIADR[21]), .D(n313), 
        .E(SIHCIADR1[21]), .F(n329), .Y(n263) );
    zao222b U226 ( .A(IHCIADR1[20]), .B(n312), .C(PERHCIADR[20]), .D(n328), 
        .E(SIHCIADR1[20]), .F(n314), .Y(n261) );
    zao222b U227 ( .A(IHCIADR1[19]), .B(n327), .C(PERHCIADR[19]), .D(n313), 
        .E(SIHCIADR1[19]), .F(n329), .Y(n259) );
    zao222b U228 ( .A(IHCIADR1[18]), .B(n312), .C(PERHCIADR[18]), .D(n328), 
        .E(SIHCIADR1[18]), .F(n314), .Y(n257) );
    zao222b U229 ( .A(IHCIADR1[17]), .B(n327), .C(PERHCIADR[17]), .D(n313), 
        .E(SIHCIADR1[17]), .F(n314), .Y(n255) );
    zao222b U230 ( .A(IHCIADR1[16]), .B(n312), .C(PERHCIADR[16]), .D(n328), 
        .E(SIHCIADR1[16]), .F(n329), .Y(n253) );
    zao222b U231 ( .A(IHCIADR1[15]), .B(n312), .C(PERHCIADR[15]), .D(n313), 
        .E(SIHCIADR1[15]), .F(n329), .Y(n251) );
    zao222b U232 ( .A(IHCIADR1[14]), .B(n327), .C(PERHCIADR[14]), .D(n328), 
        .E(SIHCIADR1[14]), .F(n314), .Y(n249) );
    zao222b U233 ( .A(IHCIADR1[13]), .B(n327), .C(PERHCIADR[13]), .D(n313), 
        .E(SIHCIADR1[13]), .F(n329), .Y(n247) );
    zao222b U234 ( .A(IHCIADR1[12]), .B(n312), .C(PERHCIADR[12]), .D(n328), 
        .E(SIHCIADR1[12]), .F(n314), .Y(n245) );
    zao222b U235 ( .A(IHCIADR1[3]), .B(n327), .C(PERHCIADR[3]), .D(n313), .E(
        SIHCIADR1[3]), .F(n329), .Y(n227) );
    zao222b U236 ( .A(IHCIADR1[2]), .B(n312), .C(PERHCIADR[2]), .D(n328), .E(
        SIHCIADR1[2]), .F(n314), .Y(n225) );
    zao222b U237 ( .A(SIHCIADD1[9]), .B(n321), .C(QHCIADD1[9]), .D(n322), .E(
        IHCIADD1[9]), .F(n323), .Y(n189) );
    zao222b U238 ( .A(SIHCIADD2[9]), .B(n324), .C(QHCIADD2[9]), .D(n325), .E(
        IHCIADD2[9]), .F(n326), .Y(n190) );
    zao222b U239 ( .A(SIHCIADD1[8]), .B(n315), .C(QHCIADD1[8]), .D(n316), .E(
        IHCIADD1[8]), .F(n317), .Y(n223) );
    zao222b U240 ( .A(SIHCIADD2[8]), .B(n318), .C(QHCIADD2[8]), .D(n319), .E(
        IHCIADD2[8]), .F(n320), .Y(n224) );
    zao222b U241 ( .A(SIHCIADD1[7]), .B(n321), .C(QHCIADD1[7]), .D(n322), .E(
        IHCIADD1[7]), .F(n323), .Y(n195) );
    zao222b U242 ( .A(SIHCIADD2[7]), .B(n324), .C(QHCIADD2[7]), .D(n325), .E(
        IHCIADD2[7]), .F(n326), .Y(n196) );
    zao222b U243 ( .A(SIHCIADD1[6]), .B(n315), .C(QHCIADD1[6]), .D(n316), .E(
        IHCIADD1[6]), .F(n317), .Y(n211) );
    zao222b U244 ( .A(SIHCIADD2[6]), .B(n318), .C(QHCIADD2[6]), .D(n319), .E(
        IHCIADD2[6]), .F(n320), .Y(n212) );
    zao222b U245 ( .A(SIHCIADD1[5]), .B(n321), .C(QHCIADD1[5]), .D(n322), .E(
        IHCIADD1[5]), .F(n323), .Y(n203) );
    zao222b U246 ( .A(SIHCIADD2[5]), .B(n324), .C(QHCIADD2[5]), .D(n325), .E(
        IHCIADD2[5]), .F(n326), .Y(n204) );
    zao222b U247 ( .A(SIHCIADD1[4]), .B(n315), .C(QHCIADD1[4]), .D(n316), .E(
        IHCIADD1[4]), .F(n317), .Y(n183) );
    zao222b U248 ( .A(SIHCIADD2[4]), .B(n318), .C(QHCIADD2[4]), .D(n319), .E(
        IHCIADD2[4]), .F(n320), .Y(n184) );
    zao222b U249 ( .A(SIHCIADD1[31]), .B(n321), .C(QHCIADD1[31]), .D(n322), 
        .E(IHCIADD1[31]), .F(n323), .Y(n167) );
    zao222b U250 ( .A(SIHCIADD2[31]), .B(n324), .C(QHCIADD2[31]), .D(n325), 
        .E(IHCIADD2[31]), .F(n326), .Y(n168) );
    zao222b U251 ( .A(SIHCIADD1[30]), .B(n315), .C(QHCIADD1[30]), .D(n316), 
        .E(IHCIADD1[30]), .F(n317), .Y(n169) );
    zao222b U252 ( .A(SIHCIADD2[30]), .B(n318), .C(QHCIADD2[30]), .D(n319), 
        .E(IHCIADD2[30]), .F(n320), .Y(n170) );
    zao222b U253 ( .A(SIHCIADD1[3]), .B(n321), .C(QHCIADD1[3]), .D(n322), .E(
        IHCIADD1[3]), .F(n323), .Y(n173) );
    zao222b U254 ( .A(SIHCIADD2[3]), .B(n324), .C(QHCIADD2[3]), .D(n325), .E(
        IHCIADD2[3]), .F(n326), .Y(n174) );
    zao222b U255 ( .A(SIHCIADD1[29]), .B(n315), .C(QHCIADD1[29]), .D(n316), 
        .E(IHCIADD1[29]), .F(n317), .Y(n179) );
    zao222b U256 ( .A(SIHCIADD2[29]), .B(n318), .C(QHCIADD2[29]), .D(n319), 
        .E(IHCIADD2[29]), .F(n320), .Y(n180) );
    zao222b U257 ( .A(SIHCIADD1[28]), .B(n321), .C(QHCIADD1[28]), .D(n322), 
        .E(IHCIADD1[28]), .F(n323), .Y(n209) );
    zao222b U258 ( .A(SIHCIADD2[28]), .B(n324), .C(QHCIADD2[28]), .D(n325), 
        .E(IHCIADD2[28]), .F(n326), .Y(n210) );
    zao222b U259 ( .A(SIHCIADD1[27]), .B(n315), .C(QHCIADD1[27]), .D(n316), 
        .E(IHCIADD1[27]), .F(n317), .Y(n197) );
    zao222b U260 ( .A(SIHCIADD2[27]), .B(n318), .C(QHCIADD2[27]), .D(n319), 
        .E(IHCIADD2[27]), .F(n320), .Y(n198) );
    zao222b U261 ( .A(SIHCIADD1[26]), .B(n321), .C(QHCIADD1[26]), .D(n322), 
        .E(IHCIADD1[26]), .F(n323), .Y(n217) );
    zao222b U262 ( .A(SIHCIADD2[26]), .B(n324), .C(QHCIADD2[26]), .D(n325), 
        .E(IHCIADD2[26]), .F(n326), .Y(n218) );
    zao222b U263 ( .A(SIHCIADD1[25]), .B(n315), .C(QHCIADD1[25]), .D(n316), 
        .E(IHCIADD1[25]), .F(n317), .Y(n193) );
    zao222b U264 ( .A(SIHCIADD2[25]), .B(n318), .C(QHCIADD2[25]), .D(n319), 
        .E(IHCIADD2[25]), .F(n320), .Y(n194) );
    zao222b U265 ( .A(SIHCIADD1[24]), .B(n321), .C(QHCIADD1[24]), .D(n322), 
        .E(IHCIADD1[24]), .F(n323), .Y(n185) );
    zao222b U266 ( .A(SIHCIADD2[24]), .B(n324), .C(QHCIADD2[24]), .D(n325), 
        .E(IHCIADD2[24]), .F(n326), .Y(n186) );
    zao222b U267 ( .A(SIHCIADD1[23]), .B(n315), .C(QHCIADD1[23]), .D(n316), 
        .E(IHCIADD1[23]), .F(n317), .Y(n161) );
    zao222b U268 ( .A(SIHCIADD2[23]), .B(n318), .C(QHCIADD2[23]), .D(n319), 
        .E(IHCIADD2[23]), .F(n320), .Y(n162) );
    zao222b U269 ( .A(SIHCIADD1[22]), .B(n321), .C(QHCIADD1[22]), .D(n322), 
        .E(IHCIADD1[22]), .F(n323), .Y(n191) );
    zao222b U270 ( .A(SIHCIADD2[22]), .B(n324), .C(QHCIADD2[22]), .D(n325), 
        .E(IHCIADD2[22]), .F(n326), .Y(n192) );
    zao222b U271 ( .A(SIHCIADD1[21]), .B(n315), .C(QHCIADD1[21]), .D(n316), 
        .E(IHCIADD1[21]), .F(n317), .Y(n221) );
    zao222b U272 ( .A(SIHCIADD2[21]), .B(n318), .C(QHCIADD2[21]), .D(n319), 
        .E(IHCIADD2[21]), .F(n320), .Y(n222) );
    zao222b U273 ( .A(SIHCIADD1[20]), .B(n321), .C(QHCIADD1[20]), .D(n322), 
        .E(IHCIADD1[20]), .F(n323), .Y(n213) );
    zao222b U274 ( .A(SIHCIADD2[20]), .B(n324), .C(QHCIADD2[20]), .D(n325), 
        .E(IHCIADD2[20]), .F(n326), .Y(n214) );
    zao222b U275 ( .A(SIHCIADD1[2]), .B(n315), .C(QHCIADD1[2]), .D(n316), .E(
        IHCIADD1[2]), .F(n317), .Y(n201) );
    zao222b U276 ( .A(SIHCIADD2[2]), .B(n318), .C(QHCIADD2[2]), .D(n319), .E(
        IHCIADD2[2]), .F(n320), .Y(n202) );
    zao222b U277 ( .A(SIHCIADD1[19]), .B(n321), .C(QHCIADD1[19]), .D(n322), 
        .E(IHCIADD1[19]), .F(n323), .Y(n205) );
    zao222b U278 ( .A(SIHCIADD2[19]), .B(n324), .C(QHCIADD2[19]), .D(n325), 
        .E(IHCIADD2[19]), .F(n326), .Y(n206) );
    zao222b U279 ( .A(SIHCIADD1[18]), .B(n315), .C(QHCIADD1[18]), .D(n316), 
        .E(IHCIADD1[18]), .F(n317), .Y(n175) );
    zao222b U280 ( .A(SIHCIADD2[18]), .B(n318), .C(QHCIADD2[18]), .D(n319), 
        .E(IHCIADD2[18]), .F(n320), .Y(n176) );
    zao222b U281 ( .A(SIHCIADD1[17]), .B(n321), .C(QHCIADD1[17]), .D(n322), 
        .E(IHCIADD1[17]), .F(n323), .Y(n181) );
    zao222b U282 ( .A(SIHCIADD2[17]), .B(n324), .C(QHCIADD2[17]), .D(n325), 
        .E(IHCIADD2[17]), .F(n326), .Y(n182) );
    zao222b U283 ( .A(SIHCIADD1[16]), .B(n315), .C(QHCIADD1[16]), .D(n316), 
        .E(IHCIADD1[16]), .F(n317), .Y(n163) );
    zao222b U284 ( .A(SIHCIADD2[16]), .B(n318), .C(QHCIADD2[16]), .D(n319), 
        .E(IHCIADD2[16]), .F(n320), .Y(n164) );
    zao222b U285 ( .A(SIHCIADD1[15]), .B(n321), .C(QHCIADD1[15]), .D(n322), 
        .E(IHCIADD1[15]), .F(n323), .Y(n187) );
    zao222b U286 ( .A(SIHCIADD2[15]), .B(n324), .C(QHCIADD2[15]), .D(n325), 
        .E(IHCIADD2[15]), .F(n326), .Y(n188) );
    zao222b U287 ( .A(SIHCIADD1[14]), .B(n315), .C(QHCIADD1[14]), .D(n316), 
        .E(IHCIADD1[14]), .F(n317), .Y(n199) );
    zao222b U288 ( .A(SIHCIADD2[14]), .B(n318), .C(QHCIADD2[14]), .D(n319), 
        .E(IHCIADD2[14]), .F(n320), .Y(n200) );
    zao222b U289 ( .A(SIHCIADD1[13]), .B(n315), .C(QHCIADD1[13]), .D(n322), 
        .E(IHCIADD1[13]), .F(n323), .Y(n207) );
    zao222b U290 ( .A(SIHCIADD2[13]), .B(n318), .C(QHCIADD2[13]), .D(n325), 
        .E(IHCIADD2[13]), .F(n326), .Y(n208) );
    zao222b U291 ( .A(SIHCIADD1[12]), .B(n321), .C(QHCIADD1[12]), .D(n316), 
        .E(IHCIADD1[12]), .F(n317), .Y(n177) );
    zao222b U292 ( .A(SIHCIADD2[12]), .B(n324), .C(QHCIADD2[12]), .D(n319), 
        .E(IHCIADD2[12]), .F(n320), .Y(n178) );
    zao222b U293 ( .A(SIHCIADD1[11]), .B(n321), .C(QHCIADD1[11]), .D(n322), 
        .E(IHCIADD1[11]), .F(n323), .Y(n171) );
    zao222b U294 ( .A(SIHCIADD2[11]), .B(n324), .C(QHCIADD2[11]), .D(n325), 
        .E(IHCIADD2[11]), .F(n326), .Y(n172) );
    zao222b U295 ( .A(SIHCIADD1[10]), .B(n315), .C(QHCIADD1[10]), .D(n316), 
        .E(IHCIADD1[10]), .F(n317), .Y(n165) );
    zao222b U296 ( .A(SIHCIADD2[10]), .B(n318), .C(QHCIADD2[10]), .D(n319), 
        .E(IHCIADD2[10]), .F(n320), .Y(n166) );
    zao222b U297 ( .A(SIHCIADD1[1]), .B(n321), .C(QHCIADD1[1]), .D(n322), .E(
        IHCIADD1[1]), .F(n323), .Y(n215) );
    zao222b U298 ( .A(SIHCIADD2[1]), .B(n324), .C(QHCIADD2[1]), .D(n325), .E(
        IHCIADD2[1]), .F(n326), .Y(n216) );
    zao222b U299 ( .A(SIHCIADD1[0]), .B(n315), .C(QHCIADD1[0]), .D(n316), .E(
        IHCIADD1[0]), .F(n317), .Y(n219) );
    zao222b U300 ( .A(SIHCIADD2[0]), .B(n318), .C(QHCIADD2[0]), .D(n319), .E(
        IHCIADD2[0]), .F(n320), .Y(n220) );
endmodule


module ITDCTL ( ITD_PARSE_GO, PARSEITDEND, ITDPARSING, ITDIDLE, FRNUM, DW0, 
    DW1, DW2, DW3, DW4, DW5, DW6, DW7, DW8, DW9, DW10, DW11, DW12, DW13, DW14, 
    DW15, GEN_PERR, PCIEND, WPR, IHCIREQ, IDWNUM, IDWOFFSET, IHCIADR, IHCIADD, 
    IHCIMWR, ITDSM, TRAN_CMD, ITD_ACT, IBUI_GO, CACHE_ADDR, CACHE_INVALID, 
    CRCERR, ACTLEN, BABBLE, PIDERR, TMOUT, RXDATA0, RXDATA1, RXDATA2, RXPID, 
    TOGMATCH, SPD, EHCI_MAC_EOT, FEMPTY, TDMAEND, IRXERR, ICMDSTART_REQ, 
    ICMDSTART, IEOT, HCI_PRESOF, LTINT_PCLK, USBINT_EN, ERRINT_EN, USBINT, 
    ERRINT, ITDIOCINT_S, ITDERRINT_S, ITDIOCINT, RECOVERYMODE, PCICLK, 
    EHCIFLOW_PCLK, TRST_ );
input  [13:0] FRNUM;
input  [31:0] DW0;
input  [31:0] DW14;
input  [31:0] DW7;
input  [31:0] DW9;
input  [7:0] RXPID;
output [3:0] IDWOFFSET;
input  [26:0] CACHE_ADDR;
input  [31:0] DW1;
input  [31:0] DW6;
input  [31:0] DW12;
input  [31:0] DW13;
output [31:0] IHCIADD;
output [31:0] IHCIADR;
input  [31:0] DW2;
input  [31:0] DW3;
input  [31:0] DW8;
input  [31:0] DW15;
input  [31:0] WPR;
input  [31:0] DW4;
input  [10:0] ACTLEN;
input  [31:0] DW5;
input  [31:0] DW10;
output [13:0] ITDSM;
input  [31:0] DW11;
output [104:0] TRAN_CMD;
output [3:0] IDWNUM;
input  ITD_PARSE_GO, GEN_PERR, PCIEND, ITD_ACT, CRCERR, BABBLE, PIDERR, TMOUT, 
    RXDATA0, RXDATA1, RXDATA2, TOGMATCH, SPD, EHCI_MAC_EOT, FEMPTY, TDMAEND, 
    ICMDSTART, HCI_PRESOF, LTINT_PCLK, USBINT_EN, ERRINT_EN, USBINT, ERRINT, 
    RECOVERYMODE, PCICLK, EHCIFLOW_PCLK, TRST_;
output PARSEITDEND, ITDPARSING, ITDIDLE, IHCIREQ, IHCIMWR, IBUI_GO, 
    CACHE_INVALID, IRXERR, ICMDSTART_REQ, IEOT, ITDIOCINT_S, ITDERRINT_S, 
    ITDIOCINT;
    wire TR_LEN931_3, TRANSOFFSET1140_7, TR_LEN_5, PG_0, TR_LEN913_2, 
        ITDSMNXT_7, HCI_PRESOF_T432, TRANSLEN813_3, SPAREO6, HCI_PRESOF_T, 
        TRANSLEN795_7, TRANSLEN_2, TRANSLEN_11, TRANSOFFSET1141_7, 
        TR_LEN931_10, TR_LEN_11, CACHE_INVALID1402, TRANSOFFSET1141_9, 
        NXTISSTSWB, TRANSLEN795_9, TRANSOFFSET_12, TRANSOFFSET1140_12, 
        SPAREO0_, ITDSMNXT_9, SPAREO8, TRANSLEN795_11, TRANSOFFSET1140_9, 
        TRANSOFFSET1141_0, TRANSLEN_5, IEOT1283, ITDERRINT_T, TRANSLEN795_0, 
        TRANSLEN813_4, TR_LEN913_5, PG_INC472, ICMDSTART_EOT1246, SPAREO1, 
        TR_LEN_2, PHASENXT_w4usbidle, TR_LEN931_4, TRANSOFFSET1140_0, 
        TRANSOFFSET1140_8, TRANSOFFSET1141_12, SPAREO9, TRANSLEN795_10, 
        TRANSLEN795_8, PHASENXT_idle, TRANSOFFSET1141_8, TR_LEN_3, TR_LEN931_5, 
        TRANSOFFSET1140_1, TRANSLEN813_5, TR_LEN913_4, SPAREO0, TRANSLEN_4, 
        TRANSLEN795_1, TRANSOFFSET1141_1, IRXERR1209, TRANSOFFSET1141_6, 
        MULT650_1, TRANSLEN795_6, MULT_0, TRANSLEN_3, TRANSLEN_10, PG_1, 
        TR_LEN913_3, ITDSMNXT_6, TRANSLEN813_2, SPAREO7, TR_LEN931_2, 
        TRANSOFFSET1140_6, TR_LEN_4, ITDIOCINT_T1439, LENGTMAX855, ACTIVE_COM, 
        ITDIOCINT_T, TR_LEN_10, TR_LEN931_11, ITDIOCINT1476, TR_LEN913_11, 
        TR_LEN_6, TR_LEN931_0, TRANSOFFSET1140_4, SPAREO5, ITDSMNXT_4, 
        TR_LEN913_1, TRANSLEN813_0, TRANSLEN_1, TRANSLEN795_4, 
        TRANSOFFSET1141_4, PARSEITDEND_PRE, TR_LEN931_9, PG_INC, ICMDSTART_EOT, 
        TRANSLEN813_9, TR_LEN913_8, TRANSLEN_8, n1016, TRANSLEN813_11, 
        TRANSOFFSET1140_11, TRANSOFFSET1141_10, TR_LEN_8, MULT612_0, 
        TRANSOFFSET1141_3, ITDERRINT_T1513, TRANSLEN795_3, TRANSLEN_6, SPAREO2, 
        TRANSLEN813_7, TR_LEN913_6, ITDSMNXT_3, TR_LEN931_7, TRANSOFFSET1140_3, 
        TR_LEN_1, TRANSOFFSET1141_11, TR_LEN_9, LENGTMAX_PRE, 
        TRANSOFFSET1140_10, TR_LEN931_6, TRANSOFFSET1140_2, TR_LEN_0, SPAREO3, 
        SPAREO1_, TRANSLEN813_6, TR_LEN913_7, ITDSMNXT_2, TRANSLEN795_2, 
        TRANSLEN_7, MULT612_1, TRANSOFFSET1141_2, TRANSOFFSET1141_5, LDPARM, 
        TRANSLEN_0, TRANSLEN795_5, SPAREO4, ITDSMNXT_5, TR_LEN913_0, 
        TRANSLEN813_1, PG_2, TR_LEN913_10, TR_LEN_7, TR_LEN931_1, 
        TRANSOFFSET1140_5, TRANSLEN813_10, TRANSLEN_9, TRANSLEN813_8, 
        TR_LEN913_9, TR_LEN931_8, n1732, n1734, n1735, n1736, n1737, n1738, 
        n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1758, n1759, 
        n1763, n1764, n1765, n1766, n1767, n1768, n1769, add_487_carry_29, 
        add_487_carry_20, add_487_carry_15, add_487_carry_8, add_487_carry_28, 
        add_487_carry_27, add_487_carry_26, add_487_carry_12, add_487_carry_6, 
        add_487_carry_14, add_487_carry_13, add_487_carry_7, add_487_carry_24, 
        add_487_carry_23, add_487_carry_21, add_487_carry_16, add_487_carry_9, 
        add_487_carry_2, add_487_carry_18, add_487_carry_25, add_487_carry_11, 
        add_487_carry_5, add_487_carry_19, add_487_carry_10, add_487_carry_4, 
        add_487_carry_22, add_487_carry_17, add_487_carry_3, n1790, n1791, 
        n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, 
        n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, 
        n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, 
        n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, 
        n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
        sub_328_carry_8, sub_328_carry_1, sub_328_B_not_10, sub_328_B_not_8, 
        sub_328_B_not_6, sub_328_B_not_1, sub_328_carry_9, sub_328_carry_7, 
        sub_328_carry_6, sub_328_B_not_7, sub_328_B_not_9, sub_328_B_not_0, 
        sub_328_carry_2, sub_328_B_not_5, sub_328_B_not_2, sub_328_carry_11, 
        sub_328_carry_10, sub_328_carry_5, sub_328_carry_4, sub_328_B_not_4, 
        sub_328_carry_3, sub_328_B_not_3, n1840, n1841, n1842, add_353_carry_8, 
        add_353_carry_1, add_353_carry_9, add_353_carry_7, add_353_carry_6, 
        add_353_carry_2, add_353_carry_11, add_353_carry_10, add_353_carry_5, 
        add_353_carry_4, add_353_carry_3, r211_carry_8, r211_carry_1, 
        r211_carry_12, r211_carry_7, r211_carry_6, r211_carry_9, r211_carry_2, 
        r211_carry_11, r211_carry_10, r211_carry_5, r211_carry_4, r211_carry_3, 
        n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
        n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
        n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
        n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
        n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
        n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
        n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
        n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
        n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
        n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
        n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
        n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
        n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
        n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
        n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
        n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
        n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
        n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
        n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
        n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
        n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
        n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
        n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2073, 
        n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
        n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, 
        n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, 
        n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, 
        n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, 
        n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, 
        n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, 
        n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, 
        n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, 
        n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, 
        n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, 
        n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, 
        n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, 
        n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, 
        n2214, n2215, n2216, _cell_414_U49_Z_10, _cell_414_U49_Z_9, 
        _cell_414_U49_Z_8, _cell_414_U49_Z_7, _cell_414_U49_Z_6, 
        _cell_414_U49_Z_5, _cell_414_U49_Z_4, _cell_414_U49_Z_3, 
        _cell_414_U49_Z_2, _cell_414_U49_Z_1, _cell_414_U49_Z_0;
    assign IDWNUM[3] = 1'b0;
    assign IDWNUM[2] = 1'b0;
    assign IDWNUM[1] = 1'b0;
    assign IDWNUM[0] = 1'b0;
    assign IDWOFFSET[3] = 1'b0;
    assign IDWOFFSET[2] = 1'b0;
    assign IDWOFFSET[1] = 1'b0;
    assign IDWOFFSET[0] = 1'b0;
    assign IHCIADR[1] = 1'b0;
    assign IHCIADR[0] = 1'b0;
    assign IHCIADD[31] = 1'b0;
    assign IHCIADD[30] = 1'b0;
    assign TRAN_CMD[51] = 1'b1;
    assign TRAN_CMD[28] = 1'b0;
    assign TRAN_CMD[27] = 1'b0;
    assign TRAN_CMD[26] = 1'b0;
    assign TRAN_CMD[25] = 1'b0;
    assign TRAN_CMD[24] = 1'b0;
    assign TRAN_CMD[23] = 1'b0;
    assign TRAN_CMD[22] = 1'b0;
    assign TRAN_CMD[21] = 1'b0;
    assign TRAN_CMD[20] = 1'b0;
    assign TRAN_CMD[19] = 1'b0;
    assign TRAN_CMD[18] = 1'b0;
    assign TRAN_CMD[17] = 1'b0;
    assign TRAN_CMD[16] = 1'b0;
    assign TRAN_CMD[15] = 1'b0;
    assign TRAN_CMD[14] = 1'b0;
    assign TRAN_CMD[13] = 1'b0;
    assign TRAN_CMD[12] = 1'b0;
    assign TRAN_CMD[11] = 1'b0;
    assign TRAN_CMD[10] = 1'b0;
    assign TRAN_CMD[7] = 1'b0;
    assign TRAN_CMD[6] = 1'b0;
    assign TRAN_CMD[5] = 1'b0;
    assign TRAN_CMD[0] = 1'b1;
    zoai21b SPARE565 ( .A(SPAREO1), .B(LDPARM), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE562 ( .A(SPAREO0), .B(NXTISSTSWB), .C(SPAREO1_), .D(
        ACTIVE_COM), .Y(SPAREO2) );
    zaoi211b SPARE563 ( .A(SPAREO4), .B(PARSEITDEND_PRE), .C(SPAREO6), .D(1'b0
        ), .Y(SPAREO8) );
    zoai21b SPARE564 ( .A(SPAREO0), .B(SPAREO8), .C(n1732), .Y(SPAREO9) );
    znr3b SPARE566 ( .A(SPAREO2), .B(LENGTMAX_PRE), .C(SPAREO0_), .Y(SPAREO4)
         );
    zdffrb SPARE561 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE568 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE560 ( .CK(PCICLK), .D(LDPARM), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE569 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb SPARE567 ( .A(SPAREO4), .Y(SPAREO5) );
    znd2b U572 ( .A(DW10[2]), .B(n1816), .Y(n1805) );
    znd2b U573 ( .A(DW10[3]), .B(n1814), .Y(n1806) );
    znd2b U574 ( .A(n1808), .B(n1807), .Y(n1834) );
    znd2b U575 ( .A(TRANSLEN_2), .B(sub_328_B_not_2), .Y(n1808) );
    znd2b U576 ( .A(TRANSLEN_1), .B(sub_328_B_not_1), .Y(n1807) );
    znr2b U577 ( .A(n1838), .B(n1836), .Y(n1837) );
    znr2b U578 ( .A(TRANSLEN_1), .B(sub_328_B_not_1), .Y(n1838) );
    znd2b U579 ( .A(TRANSLEN_0), .B(sub_328_B_not_0), .Y(n1836) );
    znd2b U580 ( .A(DW10[4]), .B(n1815), .Y(n1801) );
    znd2b U581 ( .A(DW10[5]), .B(n1812), .Y(n1802) );
    znd2b U582 ( .A(n1804), .B(n1803), .Y(n1830) );
    znd2b U583 ( .A(TRANSLEN_4), .B(sub_328_B_not_4), .Y(n1804) );
    znd2b U584 ( .A(TRANSLEN_3), .B(sub_328_B_not_3), .Y(n1803) );
    znr2b U585 ( .A(n1835), .B(n1832), .Y(n1833) );
    znr2b U586 ( .A(n1837), .B(n1834), .Y(n1835) );
    znd2b U587 ( .A(n1806), .B(n1805), .Y(n1832) );
    znd2b U588 ( .A(DW10[6]), .B(n1813), .Y(n1797) );
    znd2b U589 ( .A(DW10[7]), .B(n1810), .Y(n1798) );
    znd2b U590 ( .A(n1800), .B(n1799), .Y(n1826) );
    znd2b U591 ( .A(TRANSLEN_6), .B(sub_328_B_not_6), .Y(n1800) );
    znd2b U592 ( .A(TRANSLEN_5), .B(sub_328_B_not_5), .Y(n1799) );
    znr2b U593 ( .A(n1831), .B(n1828), .Y(n1829) );
    znr2b U594 ( .A(n1833), .B(n1830), .Y(n1831) );
    znd2b U595 ( .A(n1802), .B(n1801), .Y(n1828) );
    znd2b U596 ( .A(DW10[8]), .B(n1811), .Y(n1793) );
    znd2b U597 ( .A(DW10[9]), .B(n1809), .Y(n1794) );
    znd2b U598 ( .A(n1796), .B(n1795), .Y(n1822) );
    znd2b U599 ( .A(TRANSLEN_8), .B(sub_328_B_not_8), .Y(n1796) );
    znd2b U600 ( .A(TRANSLEN_7), .B(sub_328_B_not_7), .Y(n1795) );
    znr2b U601 ( .A(n1827), .B(n1824), .Y(n1825) );
    znr2b U602 ( .A(n1829), .B(n1826), .Y(n1827) );
    znd2b U603 ( .A(n1798), .B(n1797), .Y(n1824) );
    zao3b U604 ( .A(n2034), .B(n2037), .C(n2121), .Y(n2057) );
    zan2b U605 ( .A(n2035), .B(n2036), .Y(n2034) );
    zan2b U606 ( .A(n1869), .B(n2038), .Y(n2037) );
    zoa22b U607 ( .A(n1869), .B(n2038), .C(n2035), .D(n2036), .Y(n2055) );
    zoai21b U608 ( .A(RXDATA0), .B(n2132), .C(TOGMATCH), .Y(n2192) );
    zivb U609 ( .A(SPD), .Y(n2132) );
    znr8b U610 ( .A(RXPID[0]), .B(RXPID[1]), .C(RXPID[7]), .D(RXPID[6]), .E(
        RXPID[2]), .F(RXPID[5]), .G(RXPID[3]), .H(RXPID[4]), .Y(n2062) );
    zao22b U611 ( .A(n1734), .B(n1871), .C(n2199), .D(n2118), .Y(n2200) );
    znd2b U612 ( .A(n1792), .B(n1791), .Y(n1818) );
    znd2b U613 ( .A(TRANSLEN_9), .B(sub_328_B_not_9), .Y(n1792) );
    znd2b U614 ( .A(TRANSLEN_10), .B(sub_328_B_not_10), .Y(n1791) );
    znr2b U615 ( .A(n1823), .B(n1820), .Y(n1821) );
    znr2b U616 ( .A(n1825), .B(n1822), .Y(n1823) );
    znd2b U617 ( .A(n1794), .B(n1793), .Y(n1820) );
    znr2b U618 ( .A(n1841), .B(n1840), .Y(n1842) );
    znd2b U619 ( .A(IHCIADD[12]), .B(PG_INC), .Y(n1841) );
    zor2b U620 ( .A(ITDSM[7]), .B(n2126), .Y(n2067) );
    zan3b U621 ( .A(n2055), .B(n2056), .C(n2057), .Y(n2054) );
    zaoi2x4b U622 ( .A(n2178), .B(DW4[31]), .C(n2179), .D(DW3[31]), .E(n2180), 
        .F(DW2[31]), .G(n2181), .H(DW1[31]), .Y(n1865) );
    zor2b U623 ( .A(ITDSM[8]), .B(n2056), .Y(n2066) );
    zor2b U624 ( .A(n2118), .B(n2128), .Y(n2138) );
    zxo2b U625 ( .A(n1790), .B(MULT_0), .Y(MULT650_1) );
    zor2b U626 ( .A(MULT_0), .B(n1016), .Y(n2060) );
    zao32b U627 ( .A(n2128), .B(n2117), .C(n1734), .D(n2048), .E(n1735), .Y(
        n2190) );
    zor2b U628 ( .A(TRAN_CMD[8]), .B(n2127), .Y(n2128) );
    zivb U629 ( .A(RXDATA2), .Y(n2127) );
    zivb U630 ( .A(n2128), .Y(n2199) );
    zoa22b U631 ( .A(n1921), .B(n2050), .C(FEMPTY), .D(n2051), .Y(n2049) );
    zmux21hb U632 ( .A(TRAN_CMD[50]), .B(ACTLEN[10]), .S(TRAN_CMD[9]), .Y(
        _cell_414_U49_Z_10) );
    zmux21hb U633 ( .A(TRAN_CMD[49]), .B(ACTLEN[9]), .S(n2201), .Y(
        _cell_414_U49_Z_9) );
    zmux21hb U634 ( .A(TRAN_CMD[48]), .B(ACTLEN[8]), .S(n2201), .Y(
        _cell_414_U49_Z_8) );
    zmux21hb U635 ( .A(TRAN_CMD[47]), .B(ACTLEN[7]), .S(n2202), .Y(
        _cell_414_U49_Z_7) );
    zmux21hb U636 ( .A(TRAN_CMD[46]), .B(ACTLEN[6]), .S(n2202), .Y(
        _cell_414_U49_Z_6) );
    zmux21hb U637 ( .A(TRAN_CMD[45]), .B(ACTLEN[5]), .S(n2202), .Y(
        _cell_414_U49_Z_5) );
    zmux21hb U638 ( .A(TRAN_CMD[44]), .B(ACTLEN[4]), .S(n2202), .Y(
        _cell_414_U49_Z_4) );
    zmux21hb U639 ( .A(TRAN_CMD[43]), .B(ACTLEN[3]), .S(TRAN_CMD[9]), .Y(
        _cell_414_U49_Z_3) );
    zmux21hb U640 ( .A(TRAN_CMD[42]), .B(ACTLEN[2]), .S(n2202), .Y(
        _cell_414_U49_Z_2) );
    zmux21hb U641 ( .A(TRAN_CMD[41]), .B(ACTLEN[1]), .S(n2201), .Y(
        _cell_414_U49_Z_1) );
    zmux21hb U642 ( .A(TRAN_CMD[40]), .B(ACTLEN[0]), .S(n2201), .Y(
        _cell_414_U49_Z_0) );
    zor2b U643 ( .A(ITDSM[1]), .B(ITDSM[0]), .Y(n2084) );
    zivb U644 ( .A(n2089), .Y(n2194) );
    zor2b U645 ( .A(n1740), .B(n1738), .Y(n2198) );
    zan3b U646 ( .A(ITDSM[9]), .B(n1746), .C(IHCIADD[15]), .Y(n2061) );
    zoa22b U647 ( .A(n1852), .B(TDMAEND), .C(ITDSM[2]), .D(ITDSMNXT_3), .Y(
        n2063) );
    znr6b U648 ( .A(n1853), .B(TRAN_CMD[41]), .C(TRAN_CMD[40]), .D(TRAN_CMD
        [42]), .E(TRAN_CMD[44]), .F(TRAN_CMD[43]), .Y(n1852) );
    zmux21lb U649 ( .A(n2133), .B(n1745), .S(MULT_0), .Y(n2043) );
    zan3b U650 ( .A(n1744), .B(n1925), .C(n2053), .Y(n2133) );
    zor2b U651 ( .A(MULT_0), .B(DW11[0]), .Y(n2116) );
    znr2b U652 ( .A(n1821), .B(n1818), .Y(n1819) );
    znr2b U653 ( .A(TRANSLEN_10), .B(sub_328_B_not_10), .Y(n1817) );
    zxo2b U654 ( .A(n1840), .B(n1841), .Y(PG_1) );
    zivb U655 ( .A(PG_0), .Y(n2109) );
    zxo2b U656 ( .A(IHCIADD[12]), .B(PG_INC), .Y(PG_0) );
    zivb U657 ( .A(PG_2), .Y(n2106) );
    zxo2b U658 ( .A(IHCIADD[14]), .B(n1842), .Y(PG_2) );
    zivb U659 ( .A(PG_1), .Y(n2107) );
    zaoi2x4b U660 ( .A(DW8[16]), .B(n1854), .C(DW7[16]), .D(n2209), .E(DW6[16]
        ), .F(n2210), .G(DW5[16]), .H(n2211), .Y(n2173) );
    zaoi2x4b U661 ( .A(DW4[16]), .B(n2205), .C(DW3[16]), .D(n2206), .E(DW2[16]
        ), .F(n2207), .G(DW1[16]), .H(n2208), .Y(n2172) );
    zaoi2x4b U662 ( .A(DW8[17]), .B(n2204), .C(DW7[17]), .D(n2175), .E(DW6[17]
        ), .F(n2176), .G(DW5[17]), .H(n2177), .Y(n2170) );
    zaoi2x4b U663 ( .A(DW4[17]), .B(n2178), .C(DW3[17]), .D(n2179), .E(DW2[17]
        ), .F(n2180), .G(DW1[17]), .H(n2181), .Y(n2169) );
    zaoi2x4b U664 ( .A(DW8[18]), .B(n1854), .C(DW7[18]), .D(n2209), .E(DW6[18]
        ), .F(n2210), .G(DW5[18]), .H(n2211), .Y(n2167) );
    zaoi2x4b U665 ( .A(DW4[18]), .B(n2205), .C(DW3[18]), .D(n2206), .E(DW2[18]
        ), .F(n2207), .G(DW1[18]), .H(n2208), .Y(n2166) );
    zaoi2x4b U666 ( .A(DW8[19]), .B(n2204), .C(DW7[19]), .D(n2175), .E(DW6[19]
        ), .F(n2176), .G(DW5[19]), .H(n2177), .Y(n2164) );
    zaoi2x4b U667 ( .A(DW4[19]), .B(n2178), .C(DW3[19]), .D(n2179), .E(DW2[19]
        ), .F(n2180), .G(DW1[19]), .H(n2181), .Y(n2163) );
    zaoi2x4b U668 ( .A(DW8[20]), .B(n1854), .C(DW7[20]), .D(n2209), .E(DW6[20]
        ), .F(n2210), .G(DW5[20]), .H(n2211), .Y(n2161) );
    zaoi2x4b U669 ( .A(DW4[20]), .B(n2205), .C(DW3[20]), .D(n2206), .E(DW2[20]
        ), .F(n2207), .G(DW1[20]), .H(n2208), .Y(n2160) );
    zaoi2x4b U670 ( .A(DW8[21]), .B(n2204), .C(DW7[21]), .D(n2175), .E(DW6[21]
        ), .F(n2176), .G(DW5[21]), .H(n2177), .Y(n2158) );
    zaoi2x4b U671 ( .A(DW4[21]), .B(n2178), .C(DW3[21]), .D(n2179), .E(DW2[21]
        ), .F(n2180), .G(DW1[21]), .H(n2181), .Y(n2157) );
    zaoi2x4b U672 ( .A(DW8[22]), .B(n1854), .C(DW7[22]), .D(n2209), .E(DW6[22]
        ), .F(n2210), .G(DW5[22]), .H(n2211), .Y(n2155) );
    zaoi2x4b U673 ( .A(DW4[22]), .B(n2205), .C(DW3[22]), .D(n2206), .E(DW2[22]
        ), .F(n2207), .G(DW1[22]), .H(n2208), .Y(n2154) );
    zaoi2x4b U674 ( .A(DW8[23]), .B(n2204), .C(DW7[23]), .D(n2175), .E(DW6[23]
        ), .F(n2176), .G(DW5[23]), .H(n2177), .Y(n2152) );
    zaoi2x4b U675 ( .A(DW4[23]), .B(n2178), .C(DW3[23]), .D(n2179), .E(DW2[23]
        ), .F(n2180), .G(DW1[23]), .H(n2181), .Y(n2151) );
    zaoi2x4b U676 ( .A(DW8[24]), .B(n1854), .C(DW7[24]), .D(n2209), .E(DW6[24]
        ), .F(n2210), .G(DW5[24]), .H(n2211), .Y(n2149) );
    zaoi2x4b U677 ( .A(DW4[24]), .B(n2205), .C(DW3[24]), .D(n2206), .E(DW2[24]
        ), .F(n2207), .G(DW1[24]), .H(n2208), .Y(n2148) );
    zaoi2x4b U678 ( .A(DW8[25]), .B(n2204), .C(DW7[25]), .D(n2175), .E(DW6[25]
        ), .F(n2176), .G(DW5[25]), .H(n2177), .Y(n2146) );
    zaoi2x4b U679 ( .A(DW4[25]), .B(n2178), .C(DW3[25]), .D(n2179), .E(DW2[25]
        ), .F(n2180), .G(DW1[25]), .H(n2181), .Y(n2145) );
    zaoi2x4b U680 ( .A(DW8[26]), .B(n1854), .C(DW7[26]), .D(n2209), .E(DW6[26]
        ), .F(n2210), .G(DW5[26]), .H(n2211), .Y(n2143) );
    zaoi2x4b U681 ( .A(DW4[26]), .B(n2205), .C(DW3[26]), .D(n2206), .E(DW2[26]
        ), .F(n2207), .G(DW1[26]), .H(n2208), .Y(n2142) );
    zaoi2x4b U682 ( .A(DW8[27]), .B(n2204), .C(DW7[27]), .D(n2175), .E(DW6[27]
        ), .F(n2176), .G(DW5[27]), .H(n2177), .Y(n2140) );
    zivc U683 ( .A(n2076), .Y(n2209) );
    zivc U684 ( .A(n2077), .Y(n2210) );
    zivc U685 ( .A(n2078), .Y(n2211) );
    zaoi2x4b U686 ( .A(DW4[27]), .B(n2178), .C(DW3[27]), .D(n2179), .E(DW2[27]
        ), .F(n2180), .G(DW1[27]), .H(n2181), .Y(n2139) );
    zivc U687 ( .A(n2079), .Y(n2205) );
    zivc U688 ( .A(n2080), .Y(n2206) );
    zivc U689 ( .A(n2081), .Y(n2207) );
    zivc U690 ( .A(n2082), .Y(n2208) );
    zmux21lb U691 ( .A(n2135), .B(n2136), .S(n2137), .Y(n2134) );
    zivb U692 ( .A(n2066), .Y(n2135) );
    zivb U693 ( .A(n2067), .Y(n2137) );
    zan2b U694 ( .A(ITDSM[8]), .B(n2056), .Y(n2064) );
    zor2b U695 ( .A(ITDSM[6]), .B(ITDSM[5]), .Y(n2126) );
    zao22b U696 ( .A(ITDSM[5]), .B(ITDSM[6]), .C(n1743), .D(PCIEND), .Y(n2189)
         );
    zan2b U697 ( .A(n1925), .B(n2041), .Y(n2040) );
    zivb U698 ( .A(ACTIVE_COM), .Y(n2083) );
    znd2b U699 ( .A(n1865), .B(n1866), .Y(ACTIVE_COM) );
    zivd U700 ( .A(n1843), .Y(n2197) );
    zor2b U701 ( .A(ITDSM[3]), .B(n2070), .Y(n2071) );
    zivb U702 ( .A(PCIEND), .Y(n2124) );
    zivb U703 ( .A(n2050), .Y(n2131) );
    zivb U704 ( .A(n2060), .Y(n2088) );
    zivb U705 ( .A(n2087), .Y(n2196) );
    zmux21lb U706 ( .A(n2138), .B(n2041), .S(n1874), .Y(n1893) );
    zan2b U707 ( .A(n2190), .B(n2060), .Y(n1894) );
    zao33b U708 ( .A(n1739), .B(n1849), .C(n1850), .D(ICMDSTART), .E(n1738), 
        .F(n1851), .Y(ITDSMNXT_3) );
    zor2b U709 ( .A(IHCIADD[28]), .B(n1732), .Y(n1923) );
    zivc U710 ( .A(n2123), .Y(n1873) );
    zao22b U711 ( .A(TR_LEN913_11), .B(n1919), .C(TR_LEN_11), .D(n1736), .Y(
        TR_LEN931_11) );
    zao22b U712 ( .A(TR_LEN913_10), .B(n1919), .C(TR_LEN_10), .D(n1736), .Y(
        TR_LEN931_10) );
    zao22b U713 ( .A(n1919), .B(TR_LEN913_9), .C(n1736), .D(TR_LEN_9), .Y(
        TR_LEN931_9) );
    zao22b U714 ( .A(TR_LEN913_8), .B(n1919), .C(TR_LEN_8), .D(n1736), .Y(
        TR_LEN931_8) );
    zao22b U715 ( .A(TR_LEN913_7), .B(n1919), .C(TR_LEN_7), .D(n1736), .Y(
        TR_LEN931_7) );
    zao22b U716 ( .A(TR_LEN913_6), .B(n1919), .C(TR_LEN_6), .D(n1736), .Y(
        TR_LEN931_6) );
    zao22b U717 ( .A(TR_LEN913_5), .B(n1919), .C(TR_LEN_5), .D(n1736), .Y(
        TR_LEN931_5) );
    zao22b U718 ( .A(TR_LEN913_4), .B(n1919), .C(TR_LEN_4), .D(n1736), .Y(
        TR_LEN931_4) );
    zao22b U719 ( .A(TR_LEN913_3), .B(n1919), .C(TR_LEN_3), .D(n1736), .Y(
        TR_LEN931_3) );
    zao22b U720 ( .A(TR_LEN913_2), .B(n1919), .C(TR_LEN_2), .D(n1736), .Y(
        TR_LEN931_2) );
    zao22b U721 ( .A(TR_LEN913_1), .B(n1919), .C(TR_LEN_1), .D(n1736), .Y(
        TR_LEN931_1) );
    zao22b U722 ( .A(TR_LEN913_0), .B(n1919), .C(TR_LEN_0), .D(n1736), .Y(
        TR_LEN931_0) );
    zivc U723 ( .A(n2094), .Y(n1919) );
    zor2b U724 ( .A(IHCIADD[28]), .B(n2092), .Y(n2094) );
    zivd U725 ( .A(n2059), .Y(n1891) );
    zan2b U726 ( .A(n1862), .B(n1869), .Y(HCI_PRESOF_T432) );
    zao33b U727 ( .A(n1741), .B(n1849), .C(n1850), .D(n1740), .E(ICMDSTART), 
        .F(n1851), .Y(ITDSMNXT_5) );
    zao32b U728 ( .A(n1738), .B(n1888), .C(n1851), .D(n1889), .E(TRAN_CMD[8]), 
        .Y(ITDSMNXT_2) );
    zao32b U729 ( .A(n1740), .B(n1888), .C(n1851), .D(n1889), .E(TRAN_CMD[9]), 
        .Y(ITDSMNXT_4) );
    zivb U730 ( .A(ICMDSTART), .Y(n1888) );
    zivb U731 ( .A(n2129), .Y(n1851) );
    zor2b U732 ( .A(GEN_PERR), .B(n1862), .Y(n2129) );
    zivb U733 ( .A(n2130), .Y(n1889) );
    znd2b U734 ( .A(n1858), .B(n1859), .Y(PARSEITDEND_PRE) );
    zivb U735 ( .A(ITD_PARSE_GO), .Y(n1870) );
    zan3b U736 ( .A(n1854), .B(ITDSM[9]), .C(PHASENXT_idle), .Y(
        CACHE_INVALID1402) );
    zivb U737 ( .A(FRNUM[1]), .Y(n2073) );
    zivb U738 ( .A(FRNUM[2]), .Y(n2074) );
    zoa211b U739 ( .A(ITDIOCINT), .B(n1867), .C(n1868), .D(USBINT_EN), .Y(
        ITDIOCINT1476) );
    znd2b U740 ( .A(USBINT), .B(LTINT_PCLK), .Y(n1868) );
    zan3b U741 ( .A(n1741), .B(n1849), .C(n1890), .Y(ITDSMNXT_6) );
    zor2b U742 ( .A(ICMDSTART), .B(n1857), .Y(n1850) );
    zivb U743 ( .A(EHCI_MAC_EOT), .Y(n1857) );
    zivb U744 ( .A(n2090), .Y(PHASENXT_w4usbidle) );
    znd2b U745 ( .A(n2091), .B(n1849), .Y(n2090) );
    zor2b U746 ( .A(IHCIADD[28]), .B(BABBLE), .Y(n1921) );
    zan2b U747 ( .A(ITDERRINT_T), .B(n1920), .Y(n1922) );
    zivb U748 ( .A(n2051), .Y(n2195) );
    zivb U749 ( .A(GEN_PERR), .Y(n1849) );
    zor2b U750 ( .A(HCI_PRESOF), .B(HCI_PRESOF_T), .Y(n1862) );
    zor2b U751 ( .A(ITDSM[2]), .B(ITDSM[4]), .Y(n1863) );
    zan2b U752 ( .A(n1890), .B(ITDSM[3]), .Y(n1864) );
    zivb U753 ( .A(n1850), .Y(n1890) );
    zao21b U754 ( .A(ITDIOCINT_T), .B(n1920), .C(n1867), .Y(ITDIOCINT_T1439)
         );
    zivb U755 ( .A(LTINT_PCLK), .Y(n1920) );
    zor2b U756 ( .A(n2061), .B(GEN_PERR), .Y(n1867) );
    zmux21lb U757 ( .A(n2053), .B(n2086), .S(n1765), .Y(LENGTMAX855) );
    zivd U758 ( .A(n1858), .Y(LDPARM) );
    zor2b U759 ( .A(n1869), .B(n2090), .Y(n1858) );
    zivc U760 ( .A(n1858), .Y(n1874) );
    zan2b U761 ( .A(ITDERRINT_T), .B(LTINT_PCLK), .Y(ITDERRINT_S) );
    zan2b U762 ( .A(LTINT_PCLK), .B(ITDIOCINT_T), .Y(ITDIOCINT_S) );
    zan2b U763 ( .A(n1860), .B(n1861), .Y(ICMDSTART_REQ) );
    zivb U764 ( .A(n1924), .Y(IBUI_GO) );
    zor2b U765 ( .A(ITDSM[1]), .B(n2090), .Y(n1924) );
    zao32b U766 ( .A(n1871), .B(DW11[0]), .C(n1744), .D(n1872), .E(n2201), .Y(
        TRAN_CMD[2]) );
    zivb U767 ( .A(n2118), .Y(n1872) );
    zor2b U768 ( .A(n2048), .B(n1790), .Y(n2118) );
    zao32b U769 ( .A(n1871), .B(n1925), .C(n1744), .D(n1016), .E(n1926), .Y(
        TRAN_CMD[3]) );
    zivb U770 ( .A(n2117), .Y(n1871) );
    zor2b U771 ( .A(n1016), .B(n2048), .Y(n2117) );
    zivb U772 ( .A(DW11[0]), .Y(n1925) );
    zao21b U773 ( .A(n1745), .B(n2048), .C(TRAN_CMD[9]), .Y(n1926) );
    zmux21lb U774 ( .A(n2046), .B(n2042), .S(n1016), .Y(TRAN_CMD[4]) );
    zivb U775 ( .A(DW11[1]), .Y(n2041) );
    zivb U776 ( .A(n2116), .Y(n2047) );
    zan2b U777 ( .A(n2043), .B(n2044), .Y(n2042) );
    zivb U778 ( .A(LENGTMAX_PRE), .Y(n2053) );
    zao22b U779 ( .A(DW14[12]), .B(n2185), .C(DW13[12]), .D(n2215), .Y(n1995)
         );
    zao22b U780 ( .A(DW14[13]), .B(n2216), .C(DW13[13]), .D(n2184), .Y(n1997)
         );
    zao22b U781 ( .A(DW14[14]), .B(n2185), .C(DW13[14]), .D(n2215), .Y(n1999)
         );
    zao22b U782 ( .A(DW14[15]), .B(n2216), .C(DW13[15]), .D(n2184), .Y(n2001)
         );
    zao22b U783 ( .A(DW14[16]), .B(n2185), .C(DW13[16]), .D(n2215), .Y(n2003)
         );
    zao22b U784 ( .A(DW14[17]), .B(n2216), .C(DW13[17]), .D(n2184), .Y(n2005)
         );
    zao22b U785 ( .A(DW14[18]), .B(n2185), .C(DW13[18]), .D(n2215), .Y(n2007)
         );
    zao22b U786 ( .A(DW14[19]), .B(n2216), .C(DW13[19]), .D(n2184), .Y(n2009)
         );
    zao22b U787 ( .A(DW14[20]), .B(n2185), .C(DW13[20]), .D(n2215), .Y(n2011)
         );
    zao22b U788 ( .A(DW14[21]), .B(n2216), .C(DW13[21]), .D(n2184), .Y(n2013)
         );
    zao22b U789 ( .A(DW14[22]), .B(n2185), .C(DW13[22]), .D(n2215), .Y(n2015)
         );
    zao22b U790 ( .A(DW14[23]), .B(n2216), .C(DW13[23]), .D(n2184), .Y(n2017)
         );
    zao22b U791 ( .A(DW14[24]), .B(n2185), .C(DW13[24]), .D(n2215), .Y(n2019)
         );
    zao22b U792 ( .A(DW14[25]), .B(n2216), .C(DW13[25]), .D(n2184), .Y(n2021)
         );
    zao22b U793 ( .A(DW14[26]), .B(n2185), .C(DW13[26]), .D(n2215), .Y(n2023)
         );
    zao22b U794 ( .A(n2185), .B(DW14[27]), .C(n2215), .D(DW13[27]), .Y(n2025)
         );
    zao22b U795 ( .A(DW14[28]), .B(n2216), .C(DW13[28]), .D(n2184), .Y(n2027)
         );
    zao22b U796 ( .A(DW14[29]), .B(n2185), .C(DW13[29]), .D(n2215), .Y(n2029)
         );
    zao22b U797 ( .A(DW14[30]), .B(n2216), .C(DW13[30]), .D(n2184), .Y(n2031)
         );
    zao22b U798 ( .A(DW14[31]), .B(n2185), .C(DW13[31]), .D(n2215), .Y(n2033)
         );
    zao22b U799 ( .A(DW12[12]), .B(n2184), .C(DW13[12]), .D(n2216), .Y(n1992)
         );
    zao22b U800 ( .A(DW12[13]), .B(n2215), .C(DW13[13]), .D(n2185), .Y(n1989)
         );
    zao22b U801 ( .A(DW12[14]), .B(n2184), .C(DW13[14]), .D(n2216), .Y(n1986)
         );
    zao22b U802 ( .A(DW12[15]), .B(n2215), .C(DW13[15]), .D(n2185), .Y(n1983)
         );
    zao22b U803 ( .A(DW12[16]), .B(n2184), .C(DW13[16]), .D(n2216), .Y(n1980)
         );
    zao22b U804 ( .A(DW12[17]), .B(n2215), .C(DW13[17]), .D(n2185), .Y(n1977)
         );
    zao22b U805 ( .A(DW12[18]), .B(n2184), .C(DW13[18]), .D(n2216), .Y(n1974)
         );
    zao22b U806 ( .A(DW12[19]), .B(n2215), .C(DW13[19]), .D(n2185), .Y(n1971)
         );
    zao22b U807 ( .A(DW12[20]), .B(n2184), .C(DW13[20]), .D(n2216), .Y(n1968)
         );
    zao22b U808 ( .A(DW12[21]), .B(n2215), .C(DW13[21]), .D(n2185), .Y(n1965)
         );
    zao22b U809 ( .A(DW12[22]), .B(n2184), .C(DW13[22]), .D(n2216), .Y(n1962)
         );
    zao22b U810 ( .A(DW12[23]), .B(n2215), .C(DW13[23]), .D(n2185), .Y(n1959)
         );
    zao22b U811 ( .A(DW12[24]), .B(n2184), .C(DW13[24]), .D(n2216), .Y(n1956)
         );
    zao22b U812 ( .A(DW12[25]), .B(n2215), .C(DW13[25]), .D(n2185), .Y(n1953)
         );
    zao22b U813 ( .A(DW12[26]), .B(n2184), .C(DW13[26]), .D(n2216), .Y(n1950)
         );
    zao22b U814 ( .A(n2184), .B(DW12[27]), .C(n2216), .D(DW13[27]), .Y(n1947)
         );
    zao22b U815 ( .A(DW12[28]), .B(n2184), .C(DW13[28]), .D(n2216), .Y(n1944)
         );
    zao22b U816 ( .A(DW12[29]), .B(n2215), .C(DW13[29]), .D(n2185), .Y(n1941)
         );
    zivf U817 ( .A(n2114), .Y(n2186) );
    zivf U818 ( .A(n2113), .Y(n2187) );
    zivf U819 ( .A(n2115), .Y(n2188) );
    zao22b U820 ( .A(DW12[30]), .B(n2184), .C(DW13[30]), .D(n2216), .Y(n1938)
         );
    zivf U821 ( .A(n2112), .Y(n2184) );
    zivf U822 ( .A(n2111), .Y(n2216) );
    zivf U823 ( .A(n2110), .Y(n2182) );
    zivf U824 ( .A(n2114), .Y(n2212) );
    zivf U825 ( .A(n2113), .Y(n2213) );
    zivf U826 ( .A(n2115), .Y(n2214) );
    zao22b U827 ( .A(DW12[31]), .B(n2215), .C(DW13[31]), .D(n2185), .Y(n1935)
         );
    zivf U828 ( .A(n2112), .Y(n2215) );
    zivf U829 ( .A(n2111), .Y(n2185) );
    znd2b U830 ( .A(n1917), .B(n1918), .Y(IHCIADD[0]) );
    zaoi2x4b U831 ( .A(DW4[0]), .B(n2205), .C(DW3[0]), .D(n2206), .E(DW2[0]), 
        .F(n2207), .G(DW1[0]), .H(n2208), .Y(n1917) );
    zaoi2x4b U832 ( .A(DW8[0]), .B(n1854), .C(DW7[0]), .D(n2209), .E(DW6[0]), 
        .F(n2210), .G(DW5[0]), .H(n2211), .Y(n1918) );
    znd2b U833 ( .A(n1915), .B(n1916), .Y(IHCIADD[1]) );
    zaoi2x4b U834 ( .A(DW4[1]), .B(n2178), .C(DW3[1]), .D(n2179), .E(DW2[1]), 
        .F(n2180), .G(DW1[1]), .H(n2181), .Y(n1915) );
    zaoi2x4b U835 ( .A(DW8[1]), .B(n2204), .C(DW7[1]), .D(n2175), .E(DW6[1]), 
        .F(n2176), .G(DW5[1]), .H(n2177), .Y(n1916) );
    znd2b U836 ( .A(n1913), .B(n1914), .Y(IHCIADD[2]) );
    zaoi2x4b U837 ( .A(DW4[2]), .B(n2205), .C(DW3[2]), .D(n2206), .E(DW2[2]), 
        .F(n2207), .G(DW1[2]), .H(n2208), .Y(n1913) );
    zaoi2x4b U838 ( .A(DW8[2]), .B(n1854), .C(DW7[2]), .D(n2209), .E(DW6[2]), 
        .F(n2210), .G(DW5[2]), .H(n2211), .Y(n1914) );
    znd2b U839 ( .A(n1911), .B(n1912), .Y(IHCIADD[3]) );
    zaoi2x4b U840 ( .A(DW4[3]), .B(n2178), .C(DW3[3]), .D(n2179), .E(DW2[3]), 
        .F(n2180), .G(DW1[3]), .H(n2181), .Y(n1911) );
    zaoi2x4b U841 ( .A(DW8[3]), .B(n2204), .C(DW7[3]), .D(n2175), .E(DW6[3]), 
        .F(n2176), .G(DW5[3]), .H(n2177), .Y(n1912) );
    znd2b U842 ( .A(n1909), .B(n1910), .Y(IHCIADD[4]) );
    zaoi2x4b U843 ( .A(DW4[4]), .B(n2205), .C(DW3[4]), .D(n2206), .E(DW2[4]), 
        .F(n2207), .G(DW1[4]), .H(n2208), .Y(n1909) );
    zaoi2x4b U844 ( .A(DW8[4]), .B(n1854), .C(DW7[4]), .D(n2209), .E(DW6[4]), 
        .F(n2210), .G(DW5[4]), .H(n2211), .Y(n1910) );
    znd2b U845 ( .A(n1907), .B(n1908), .Y(IHCIADD[5]) );
    zaoi2x4b U846 ( .A(DW4[5]), .B(n2178), .C(DW3[5]), .D(n2179), .E(DW2[5]), 
        .F(n2180), .G(DW1[5]), .H(n2181), .Y(n1907) );
    zaoi2x4b U847 ( .A(DW8[5]), .B(n2204), .C(DW7[5]), .D(n2175), .E(DW6[5]), 
        .F(n2176), .G(DW5[5]), .H(n2177), .Y(n1908) );
    znd2b U848 ( .A(n1905), .B(n1906), .Y(IHCIADD[6]) );
    zaoi2x4b U849 ( .A(DW4[6]), .B(n2205), .C(DW3[6]), .D(n2206), .E(DW2[6]), 
        .F(n2207), .G(DW1[6]), .H(n2208), .Y(n1905) );
    zaoi2x4b U850 ( .A(DW8[6]), .B(n1854), .C(DW7[6]), .D(n2209), .E(DW6[6]), 
        .F(n2210), .G(DW5[6]), .H(n2211), .Y(n1906) );
    znd2b U851 ( .A(n1903), .B(n1904), .Y(IHCIADD[7]) );
    zaoi2x4b U852 ( .A(DW4[7]), .B(n2178), .C(DW3[7]), .D(n2179), .E(DW2[7]), 
        .F(n2180), .G(DW1[7]), .H(n2181), .Y(n1903) );
    zaoi2x4b U853 ( .A(DW8[7]), .B(n2204), .C(DW7[7]), .D(n2175), .E(DW6[7]), 
        .F(n2176), .G(DW5[7]), .H(n2177), .Y(n1904) );
    znd2b U854 ( .A(n1901), .B(n1902), .Y(IHCIADD[8]) );
    zaoi2x4b U855 ( .A(DW4[8]), .B(n2205), .C(DW3[8]), .D(n2206), .E(DW2[8]), 
        .F(n2207), .G(DW1[8]), .H(n2208), .Y(n1901) );
    zaoi2x4b U856 ( .A(DW8[8]), .B(n1854), .C(DW7[8]), .D(n2209), .E(DW6[8]), 
        .F(n2210), .G(DW5[8]), .H(n2211), .Y(n1902) );
    znd2b U857 ( .A(n1899), .B(n1900), .Y(IHCIADD[9]) );
    zaoi2x4b U858 ( .A(DW4[9]), .B(n2178), .C(DW3[9]), .D(n2179), .E(DW2[9]), 
        .F(n2180), .G(DW1[9]), .H(n2181), .Y(n1899) );
    zaoi2x4b U859 ( .A(DW8[9]), .B(n2204), .C(DW7[9]), .D(n2175), .E(DW6[9]), 
        .F(n2176), .G(DW5[9]), .H(n2177), .Y(n1900) );
    znd2b U860 ( .A(n1897), .B(n1898), .Y(IHCIADD[10]) );
    zaoi2x4b U861 ( .A(DW4[10]), .B(n2205), .C(DW3[10]), .D(n2206), .E(DW2[10]
        ), .F(n2207), .G(DW1[10]), .H(n2208), .Y(n1897) );
    zaoi2x4b U862 ( .A(DW8[10]), .B(n1854), .C(DW7[10]), .D(n2209), .E(DW6[10]
        ), .F(n2210), .G(DW5[10]), .H(n2211), .Y(n1898) );
    znd2b U863 ( .A(n1895), .B(n1896), .Y(IHCIADD[11]) );
    zaoi2x4b U864 ( .A(DW4[11]), .B(n2178), .C(DW3[11]), .D(n2179), .E(DW2[11]
        ), .F(n2180), .G(DW1[11]), .H(n2181), .Y(n1895) );
    zaoi2x4b U865 ( .A(DW8[11]), .B(n2204), .C(DW7[11]), .D(n2175), .E(DW6[11]
        ), .F(n2176), .G(DW5[11]), .H(n2177), .Y(n1896) );
    znd2b U866 ( .A(n1927), .B(n1928), .Y(IHCIADD[12]) );
    zaoi2x4b U867 ( .A(DW4[12]), .B(n2205), .C(DW3[12]), .D(n2206), .E(DW2[12]
        ), .F(n2207), .G(DW1[12]), .H(n2208), .Y(n1927) );
    zaoi2x4b U868 ( .A(DW8[12]), .B(n1854), .C(DW7[12]), .D(n2209), .E(DW6[12]
        ), .F(n2210), .G(DW5[12]), .H(n2211), .Y(n1928) );
    znd2b U869 ( .A(n1929), .B(n1930), .Y(IHCIADD[13]) );
    zaoi2x4b U870 ( .A(DW4[13]), .B(n2178), .C(DW3[13]), .D(n2179), .E(DW2[13]
        ), .F(n2180), .G(DW1[13]), .H(n2181), .Y(n1929) );
    zaoi2x4b U871 ( .A(DW8[13]), .B(n2204), .C(DW7[13]), .D(n2175), .E(DW6[13]
        ), .F(n2176), .G(DW5[13]), .H(n2177), .Y(n1930) );
    zivb U872 ( .A(IHCIADD[13]), .Y(n1840) );
    znd2b U873 ( .A(n1931), .B(n1932), .Y(IHCIADD[14]) );
    zaoi2x4b U874 ( .A(DW4[14]), .B(n2205), .C(DW3[14]), .D(n2206), .E(DW2[14]
        ), .F(n2207), .G(DW1[14]), .H(n2208), .Y(n1931) );
    zaoi2x4b U875 ( .A(DW8[14]), .B(n1854), .C(DW7[14]), .D(n2209), .E(DW6[14]
        ), .F(n2210), .G(DW5[14]), .H(n2211), .Y(n1932) );
    zivd U876 ( .A(n2075), .Y(n1854) );
    znd2b U877 ( .A(n1847), .B(n1848), .Y(IHCIADD[15]) );
    zaoi2x4b U878 ( .A(DW4[15]), .B(n2178), .C(DW3[15]), .D(n2179), .E(DW2[15]
        ), .F(n2180), .G(DW1[15]), .H(n2181), .Y(n1847) );
    zivd U879 ( .A(n2079), .Y(n2178) );
    zivd U880 ( .A(n2080), .Y(n2179) );
    zivd U881 ( .A(n2081), .Y(n2180) );
    zivd U882 ( .A(n2082), .Y(n2181) );
    zaoi2x4b U883 ( .A(DW8[15]), .B(n2204), .C(DW7[15]), .D(n2175), .E(DW6[15]
        ), .F(n2176), .G(DW5[15]), .H(n2177), .Y(n1848) );
    zivd U884 ( .A(n2075), .Y(n2204) );
    zivd U885 ( .A(n2076), .Y(n2175) );
    zivd U886 ( .A(n2077), .Y(n2176) );
    zivd U887 ( .A(n2078), .Y(n2177) );
    zmux21lb U888 ( .A(n2174), .B(n2105), .S(n2201), .Y(IHCIADD[16]) );
    zivb U889 ( .A(n1887), .Y(n2174) );
    znd2b U890 ( .A(n2172), .B(n2173), .Y(n1887) );
    zmux21lb U891 ( .A(n2171), .B(n2104), .S(TRAN_CMD[9]), .Y(IHCIADD[17]) );
    zivb U892 ( .A(n1886), .Y(n2171) );
    znd2b U893 ( .A(n2169), .B(n2170), .Y(n1886) );
    zmux21lb U894 ( .A(n2168), .B(n2101), .S(n2201), .Y(IHCIADD[18]) );
    zivb U895 ( .A(n1885), .Y(n2168) );
    znd2b U896 ( .A(n2166), .B(n2167), .Y(n1885) );
    zmux21lb U897 ( .A(n2165), .B(n2100), .S(TRAN_CMD[9]), .Y(IHCIADD[19]) );
    zivb U898 ( .A(n1884), .Y(n2165) );
    znd2b U899 ( .A(n2163), .B(n2164), .Y(n1884) );
    zmux21lb U900 ( .A(n2162), .B(n2099), .S(n2201), .Y(IHCIADD[20]) );
    zivb U901 ( .A(n1883), .Y(n2162) );
    znd2b U902 ( .A(n2160), .B(n2161), .Y(n1883) );
    zmux21lb U903 ( .A(n2159), .B(n2098), .S(TRAN_CMD[9]), .Y(IHCIADD[21]) );
    zivb U904 ( .A(n1882), .Y(n2159) );
    znd2b U905 ( .A(n2157), .B(n2158), .Y(n1882) );
    zmux21lb U906 ( .A(n2156), .B(n2097), .S(n2201), .Y(IHCIADD[22]) );
    zivb U907 ( .A(n1881), .Y(n2156) );
    znd2b U908 ( .A(n2154), .B(n2155), .Y(n1881) );
    zmux21lb U909 ( .A(n2153), .B(n2096), .S(TRAN_CMD[9]), .Y(IHCIADD[23]) );
    zivb U910 ( .A(n1880), .Y(n2153) );
    znd2b U911 ( .A(n2151), .B(n2152), .Y(n1880) );
    zmux21lb U912 ( .A(n2150), .B(n2095), .S(n2201), .Y(IHCIADD[24]) );
    zivb U913 ( .A(n1879), .Y(n2150) );
    znd2b U914 ( .A(n2148), .B(n2149), .Y(n1879) );
    zmux21lb U915 ( .A(n2147), .B(n2093), .S(n2201), .Y(IHCIADD[25]) );
    zivb U916 ( .A(n1878), .Y(n2147) );
    znd2b U917 ( .A(n2145), .B(n2146), .Y(n1878) );
    zmux21lb U918 ( .A(n2144), .B(n2103), .S(n2201), .Y(IHCIADD[26]) );
    zivb U919 ( .A(n1877), .Y(n2144) );
    znd2b U920 ( .A(n2142), .B(n2143), .Y(n1877) );
    zmux21lb U921 ( .A(n2141), .B(n2102), .S(n2201), .Y(IHCIADD[27]) );
    zivb U922 ( .A(n1875), .Y(n2141) );
    znd2b U923 ( .A(n2139), .B(n2140), .Y(n1875) );
    zan2b U924 ( .A(n1855), .B(n1856), .Y(ITDPARSING) );
    zor2b U925 ( .A(GEN_PERR), .B(n1746), .Y(n1855) );
    zivb U926 ( .A(PHASENXT_idle), .Y(n1856) );
    zivb U927 ( .A(n1855), .Y(ITDSMNXT_9) );
    zdffrb TRANSLEN_reg_11 ( .CK(PCICLK), .D(TRANSLEN813_11), .R(TRST_), .Q(
        TRANSLEN_11), .QN(n1839) );
    zdffqrb TRANSLEN_reg_10 ( .CK(PCICLK), .D(TRANSLEN813_10), .R(TRST_), .Q(
        TRANSLEN_10) );
    zdffqrb TRANSLEN_reg_9 ( .CK(PCICLK), .D(TRANSLEN813_9), .R(TRST_), .Q(
        TRANSLEN_9) );
    zivb U928 ( .A(TRANSLEN_9), .Y(n1809) );
    zdffqrb TRANSLEN_reg_8 ( .CK(PCICLK), .D(TRANSLEN813_8), .R(TRST_), .Q(
        TRANSLEN_8) );
    zivb U929 ( .A(TRANSLEN_8), .Y(n1811) );
    zdffqrb TRANSLEN_reg_7 ( .CK(PCICLK), .D(TRANSLEN813_7), .R(TRST_), .Q(
        TRANSLEN_7) );
    zivb U930 ( .A(TRANSLEN_7), .Y(n1810) );
    zdffqrb TRANSLEN_reg_6 ( .CK(PCICLK), .D(TRANSLEN813_6), .R(TRST_), .Q(
        TRANSLEN_6) );
    zivb U931 ( .A(TRANSLEN_6), .Y(n1813) );
    zdffqrb TRANSLEN_reg_5 ( .CK(PCICLK), .D(TRANSLEN813_5), .R(TRST_), .Q(
        TRANSLEN_5) );
    zivb U932 ( .A(TRANSLEN_5), .Y(n1812) );
    zdffqrb TRANSLEN_reg_4 ( .CK(PCICLK), .D(TRANSLEN813_4), .R(TRST_), .Q(
        TRANSLEN_4) );
    zivb U933 ( .A(TRANSLEN_4), .Y(n1815) );
    zdffqrb TRANSLEN_reg_3 ( .CK(PCICLK), .D(TRANSLEN813_3), .R(TRST_), .Q(
        TRANSLEN_3) );
    zivb U934 ( .A(TRANSLEN_3), .Y(n1814) );
    zdffqrb TRANSLEN_reg_2 ( .CK(PCICLK), .D(TRANSLEN813_2), .R(TRST_), .Q(
        TRANSLEN_2) );
    zivb U935 ( .A(TRANSLEN_2), .Y(n1816) );
    zdffqrb TRANSLEN_reg_1 ( .CK(PCICLK), .D(TRANSLEN813_1), .R(TRST_), .Q(
        TRANSLEN_1) );
    zdffqrb TRANSLEN_reg_0 ( .CK(PCICLK), .D(TRANSLEN813_0), .R(TRST_), .Q(
        TRANSLEN_0) );
    zdffqrb TR_LEN_reg_11 ( .CK(PCICLK), .D(TR_LEN931_11), .R(TRST_), .Q(
        TR_LEN_11) );
    zivb U936 ( .A(TR_LEN_11), .Y(n2102) );
    zdffqrb TR_LEN_reg_10 ( .CK(PCICLK), .D(TR_LEN931_10), .R(TRST_), .Q(
        TR_LEN_10) );
    zivb U937 ( .A(TR_LEN_10), .Y(n2103) );
    zdffqrb TR_LEN_reg_9 ( .CK(PCICLK), .D(TR_LEN931_9), .R(TRST_), .Q(
        TR_LEN_9) );
    zivb U938 ( .A(TR_LEN_9), .Y(n2093) );
    zdffqrb TR_LEN_reg_8 ( .CK(PCICLK), .D(TR_LEN931_8), .R(TRST_), .Q(
        TR_LEN_8) );
    zivb U939 ( .A(TR_LEN_8), .Y(n2095) );
    zdffqrb TR_LEN_reg_7 ( .CK(PCICLK), .D(TR_LEN931_7), .R(TRST_), .Q(
        TR_LEN_7) );
    zivb U940 ( .A(TR_LEN_7), .Y(n2096) );
    zdffqrb TR_LEN_reg_6 ( .CK(PCICLK), .D(TR_LEN931_6), .R(TRST_), .Q(
        TR_LEN_6) );
    zivb U941 ( .A(TR_LEN_6), .Y(n2097) );
    zdffqrb TR_LEN_reg_5 ( .CK(PCICLK), .D(TR_LEN931_5), .R(TRST_), .Q(
        TR_LEN_5) );
    zivb U942 ( .A(TR_LEN_5), .Y(n2098) );
    zdffqrb TR_LEN_reg_4 ( .CK(PCICLK), .D(TR_LEN931_4), .R(TRST_), .Q(
        TR_LEN_4) );
    zivb U943 ( .A(TR_LEN_4), .Y(n2099) );
    zdffqrb TR_LEN_reg_3 ( .CK(PCICLK), .D(TR_LEN931_3), .R(TRST_), .Q(
        TR_LEN_3) );
    zivb U944 ( .A(TR_LEN_3), .Y(n2100) );
    zdffqrb TR_LEN_reg_2 ( .CK(PCICLK), .D(TR_LEN931_2), .R(TRST_), .Q(
        TR_LEN_2) );
    zivb U945 ( .A(TR_LEN_2), .Y(n2101) );
    zdffqrb TR_LEN_reg_1 ( .CK(PCICLK), .D(TR_LEN931_1), .R(TRST_), .Q(
        TR_LEN_1) );
    zivb U946 ( .A(TR_LEN_1), .Y(n2104) );
    zdffqrb TR_LEN_reg_0 ( .CK(PCICLK), .D(TR_LEN931_0), .R(TRST_), .Q(
        TR_LEN_0) );
    zivb U947 ( .A(TR_LEN_0), .Y(n2105) );
    zdffqrb TRANSOFFSET_reg_12 ( .CK(PCICLK), .D(TRANSOFFSET1140_12), .R(TRST_
        ), .Q(TRANSOFFSET_12) );
    zdffqrb TRANSOFFSET_reg_11 ( .CK(PCICLK), .D(TRANSOFFSET1140_11), .R(TRST_
        ), .Q(TRAN_CMD[83]) );
    zdffqrb TRANSOFFSET_reg_10 ( .CK(PCICLK), .D(TRANSOFFSET1140_10), .R(TRST_
        ), .Q(TRAN_CMD[82]) );
    zdffqrb TRANSOFFSET_reg_9 ( .CK(PCICLK), .D(TRANSOFFSET1140_9), .R(TRST_), 
        .Q(TRAN_CMD[81]) );
    zdffqrb TRANSOFFSET_reg_8 ( .CK(PCICLK), .D(TRANSOFFSET1140_8), .R(TRST_), 
        .Q(TRAN_CMD[80]) );
    zdffqrb TRANSOFFSET_reg_7 ( .CK(PCICLK), .D(TRANSOFFSET1140_7), .R(TRST_), 
        .Q(TRAN_CMD[79]) );
    zdffqrb TRANSOFFSET_reg_6 ( .CK(PCICLK), .D(TRANSOFFSET1140_6), .R(TRST_), 
        .Q(TRAN_CMD[78]) );
    zdffqrb TRANSOFFSET_reg_5 ( .CK(PCICLK), .D(TRANSOFFSET1140_5), .R(TRST_), 
        .Q(TRAN_CMD[77]) );
    zdffqrb TRANSOFFSET_reg_4 ( .CK(PCICLK), .D(TRANSOFFSET1140_4), .R(TRST_), 
        .Q(TRAN_CMD[76]) );
    zdffqrb TRANSOFFSET_reg_3 ( .CK(PCICLK), .D(TRANSOFFSET1140_3), .R(TRST_), 
        .Q(TRAN_CMD[75]) );
    zdffqrb TRANSOFFSET_reg_2 ( .CK(PCICLK), .D(TRANSOFFSET1140_2), .R(TRST_), 
        .Q(TRAN_CMD[74]) );
    zdffqrb TRANSOFFSET_reg_1 ( .CK(PCICLK), .D(TRANSOFFSET1140_1), .R(TRST_), 
        .Q(TRAN_CMD[73]) );
    zdffqrb TRANSOFFSET_reg_0 ( .CK(PCICLK), .D(TRANSOFFSET1140_0), .R(TRST_), 
        .Q(TRAN_CMD[72]) );
    zdffqrb HCI_PRESOF_T_reg ( .CK(PCICLK), .D(HCI_PRESOF_T432), .R(TRST_), 
        .Q(HCI_PRESOF_T) );
    zdffqrb ITDSM_reg_5 ( .CK(PCICLK), .D(ITDSMNXT_5), .R(TRST_), .Q(ITDSM[5])
         );
    zivb U948 ( .A(ITDSM[5]), .Y(n2125) );
    zdffqrb ITDSM_reg_2 ( .CK(PCICLK), .D(ITDSMNXT_2), .R(TRST_), .Q(ITDSM[2])
         );
    zivb U949 ( .A(ITDSM[2]), .Y(n2036) );
    zdffqrb PG_INC_reg ( .CK(PCICLK), .D(PG_INC472), .R(TRST_), .Q(PG_INC) );
    zdffqrb ITDSM_reg_4 ( .CK(PCICLK), .D(ITDSMNXT_4), .R(TRST_), .Q(ITDSM[4])
         );
    zivb U950 ( .A(ITDSM[4]), .Y(n2035) );
    zdffqrb ICMDSTART_EOT_reg ( .CK(PCICLK), .D(ICMDSTART_EOT1246), .R(TRST_), 
        .Q(ICMDSTART_EOT) );
    zivb U951 ( .A(ICMDSTART_EOT), .Y(n1861) );
    zdffqrb PARSEITDEND_reg ( .CK(PCICLK), .D(PARSEITDEND_PRE), .R(TRST_), .Q(
        PARSEITDEND) );
    zdffqrb CACHE_INVALID_reg ( .CK(PCICLK), .D(CACHE_INVALID1402), .R(TRST_), 
        .Q(CACHE_INVALID) );
    zdffqrb ITDIOCINT_reg ( .CK(EHCIFLOW_PCLK), .D(ITDIOCINT1476), .R(TRST_), 
        .Q(ITDIOCINT) );
    zdffqrb ITDSM_reg_6 ( .CK(PCICLK), .D(ITDSMNXT_6), .R(TRST_), .Q(ITDSM[6])
         );
    zivb U952 ( .A(ITDSM[6]), .Y(n2092) );
    zdffqrb ITDSM_reg_1 ( .CK(PCICLK), .D(PHASENXT_w4usbidle), .R(TRST_), .Q(
        ITDSM[1]) );
    zivb U953 ( .A(ITDSM[1]), .Y(n2038) );
    zdffqrb ITDERRINT_T_reg ( .CK(EHCIFLOW_PCLK), .D(ITDERRINT_T1513), .R(
        TRST_), .Q(ITDERRINT_T) );
    zdffqrb ITDSM_reg_8 ( .CK(PCICLK), .D(n1763), .R(TRST_), .Q(ITDSM[8]) );
    zivb U954 ( .A(ITDSM[8]), .Y(n2085) );
    zdffqrb IEOT_reg ( .CK(PCICLK), .D(IEOT1283), .R(TRST_), .Q(IEOT) );
    zdffqrb ITDIOCINT_T_reg ( .CK(EHCIFLOW_PCLK), .D(ITDIOCINT_T1439), .R(
        TRST_), .Q(ITDIOCINT_T) );
    zdffrb LENGTMAX_reg ( .CK(PCICLK), .D(LENGTMAX855), .R(TRST_), .QN(n2086)
         );
    zdffrb MULT_reg_1 ( .CK(PCICLK), .D(MULT612_1), .R(TRST_), .Q(n1016), .QN(
        n1790) );
    zan4b U955 ( .A(ITD_ACT), .B(ITDSM[5]), .C(EHCI_MAC_EOT), .D(n2193), .Y(
        n1732) );
    znr2b U956 ( .A(n2201), .B(n2053), .Y(TRAN_CMD[1]) );
    zan2b U957 ( .A(RXDATA1), .B(n2202), .Y(n1734) );
    znr2b U958 ( .A(n1734), .B(n2058), .Y(n1735) );
    zoa21d U959 ( .A(IHCIADD[28]), .B(n2092), .C(n1858), .Y(n1736) );
    znr4b U960 ( .A(ITDSM[1]), .B(n1863), .C(n1869), .D(n2071), .Y(n1737) );
    znr4b U961 ( .A(n2084), .B(n2036), .C(ITDSM[4]), .D(n2071), .Y(n1738) );
    znr4b U962 ( .A(n2084), .B(n2121), .C(n1863), .D(n2070), .Y(n1739) );
    znr4b U963 ( .A(n2084), .B(n2035), .C(ITDSM[2]), .D(n2071), .Y(n1740) );
    znr4b U964 ( .A(ITDSM[9]), .B(ITDSM[7]), .C(n2125), .D(n2119), .Y(n1741)
         );
    znr4b U965 ( .A(ITDSM[6]), .B(n2069), .C(n2085), .D(n2056), .Y(n1742) );
    znr4b U966 ( .A(ITDSM[7]), .B(ITDSM[5]), .C(n1759), .D(n2119), .Y(n1743)
         );
    znr2b U967 ( .A(n2201), .B(n2041), .Y(n1744) );
    znr3b U968 ( .A(n2041), .B(n1925), .C(TRAN_CMD[1]), .Y(n1745) );
    zaoi222b U969 ( .A(n1743), .B(n2124), .C(n2131), .D(n1921), .E(n1742), .F(
        n2087), .Y(n1746) );
    zmux21hb U970 ( .A(TRANSLEN_10), .B(DW10[10]), .S(LENGTMAX_PRE), .Y(
        TRAN_CMD[50]) );
    zmux21hb U971 ( .A(TRANSLEN_9), .B(DW10[9]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [49]) );
    zmux21hb U972 ( .A(TRANSLEN_8), .B(DW10[8]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [48]) );
    zmux21hb U973 ( .A(TRANSLEN_7), .B(DW10[7]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [47]) );
    zmux21hb U974 ( .A(TRANSLEN_6), .B(DW10[6]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [46]) );
    zmux21hb U975 ( .A(TRANSLEN_5), .B(DW10[5]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [45]) );
    zmux21hb U976 ( .A(TRANSLEN_4), .B(DW10[4]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [44]) );
    zmux21hb U977 ( .A(TRANSLEN_3), .B(DW10[3]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [43]) );
    zmux21hb U978 ( .A(TRANSLEN_2), .B(DW10[2]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [42]) );
    zmux21hb U979 ( .A(TRANSLEN_1), .B(DW10[1]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [41]) );
    zmux21hb U980 ( .A(TRANSLEN_0), .B(DW10[0]), .S(LENGTMAX_PRE), .Y(TRAN_CMD
        [40]) );
    zivb U981 ( .A(DW10[8]), .Y(sub_328_B_not_8) );
    zivb U982 ( .A(DW10[6]), .Y(sub_328_B_not_6) );
    zivb U983 ( .A(DW10[4]), .Y(sub_328_B_not_4) );
    zivb U984 ( .A(DW10[2]), .Y(sub_328_B_not_2) );
    zivb U985 ( .A(DW10[1]), .Y(sub_328_B_not_1) );
    zivb U986 ( .A(DW10[3]), .Y(sub_328_B_not_3) );
    zivb U987 ( .A(DW10[5]), .Y(sub_328_B_not_5) );
    zivb U988 ( .A(DW10[7]), .Y(sub_328_B_not_7) );
    zivb U989 ( .A(DW10[9]), .Y(sub_328_B_not_9) );
    zivb U990 ( .A(DW10[10]), .Y(sub_328_B_not_10) );
    zivb U991 ( .A(DW10[0]), .Y(sub_328_B_not_0) );
    zdffqrb MULT_reg_0 ( .CK(PCICLK), .D(MULT612_0), .R(TRST_), .Q(MULT_0) );
    zivb U992 ( .A(MULT_0), .Y(n2048) );
    zor2b U993 ( .A(n1819), .B(n1817), .Y(n1758) );
    zivd U994 ( .A(n2203), .Y(n2201) );
    ziv11d U995 ( .A(n2202), .Y(TRAN_CMD[8]), .Z(TRAN_CMD[9]) );
    zivb U996 ( .A(FRNUM[0]), .Y(IHCIADR[2]) );
    ziv11b U997 ( .A(ITDSM[9]), .Y(n1759), .Z(IHCIMWR) );
    zdffqrb ITDSM_reg_9 ( .CK(PCICLK), .D(ITDSMNXT_9), .R(TRST_), .Q(ITDSM[9])
         );
    zivb U998 ( .A(n2203), .Y(n2202) );
    zivb U999 ( .A(DW10[11]), .Y(n2203) );
    zdffqrb ITDSM_reg_7 ( .CK(PCICLK), .D(ITDSMNXT_7), .R(TRST_), .Q(ITDSM[7])
         );
    zor2b U1000 ( .A(GEN_PERR), .B(n2049), .Y(n2120) );
    zivb U1001 ( .A(ITDSM[3]), .Y(n2121) );
    zan2b U1002 ( .A(n2122), .B(n1849), .Y(n1763) );
    zivb U1003 ( .A(n2108), .Y(n1764) );
    zao22b U1004 ( .A(DW14[25]), .B(n2182), .C(DW15[25]), .D(n1764), .Y(n1951)
         );
    zao22b U1005 ( .A(DW14[12]), .B(n2182), .C(DW15[12]), .D(n2183), .Y(n1990)
         );
    zao22b U1006 ( .A(DW14[23]), .B(n2182), .C(DW15[23]), .D(n2183), .Y(n1957)
         );
    zao22b U1007 ( .A(DW14[26]), .B(n2182), .C(DW15[26]), .D(n2183), .Y(n1948)
         );
    zao22b U1008 ( .A(DW14[16]), .B(n2182), .C(DW15[16]), .D(n1764), .Y(n1978)
         );
    zao22b U1009 ( .A(DW14[22]), .B(n2182), .C(DW15[22]), .D(n2183), .Y(n1960)
         );
    zao22b U1010 ( .A(DW14[28]), .B(n2182), .C(DW15[28]), .D(n2183), .Y(n1942)
         );
    zao22b U1011 ( .A(DW14[14]), .B(n2182), .C(DW15[14]), .D(n2183), .Y(n1984)
         );
    zao22b U1012 ( .A(DW14[29]), .B(n2182), .C(DW15[29]), .D(n2183), .Y(n1939)
         );
    zao22b U1013 ( .A(DW14[17]), .B(n2182), .C(DW15[17]), .D(n2183), .Y(n1975)
         );
    zao22b U1014 ( .A(DW14[30]), .B(n2182), .C(DW15[30]), .D(n2183), .Y(n1936)
         );
    zao22b U1015 ( .A(DW14[24]), .B(n2182), .C(DW15[24]), .D(n2183), .Y(n1954)
         );
    zao22b U1016 ( .A(DW14[31]), .B(n2182), .C(DW15[31]), .D(n1764), .Y(n1933)
         );
    zao22b U1017 ( .A(DW14[27]), .B(n2182), .C(DW15[27]), .D(n2183), .Y(n1945)
         );
    zao22b U1018 ( .A(DW14[18]), .B(n2182), .C(DW15[18]), .D(n2183), .Y(n1972)
         );
    zao22b U1019 ( .A(DW14[13]), .B(n2182), .C(DW15[13]), .D(n1764), .Y(n1987)
         );
    zao22b U1020 ( .A(DW14[19]), .B(n2182), .C(DW15[19]), .D(n1764), .Y(n1969)
         );
    zao22b U1021 ( .A(DW14[15]), .B(n2182), .C(DW15[15]), .D(n1764), .Y(n1981)
         );
    zao22b U1022 ( .A(DW14[20]), .B(n2182), .C(DW15[20]), .D(n2183), .Y(n1966)
         );
    zao22b U1023 ( .A(DW14[21]), .B(n2182), .C(DW15[21]), .D(n1764), .Y(n1963)
         );
    zor2b U1024 ( .A(n2106), .B(n2107), .Y(n2108) );
    zivc U1025 ( .A(n2108), .Y(n2183) );
    zivd U1026 ( .A(n1765), .Y(NXTISSTSWB) );
    zivb U1027 ( .A(n1763), .Y(n1766) );
    znr2b U1028 ( .A(ITDSM[7]), .B(n2120), .Y(n1767) );
    znr2b U1029 ( .A(n2121), .B(n1766), .Y(n1768) );
    znr2b U1030 ( .A(n1767), .B(n1768), .Y(n1765) );
    zao22b U1031 ( .A(TRANSOFFSET_12), .B(n1891), .C(TRANSOFFSET1141_12), .D(
        NXTISSTSWB), .Y(TRANSOFFSET1140_12) );
    zor2b U1032 ( .A(NXTISSTSWB), .B(LDPARM), .Y(n2059) );
    zdffqrb ITDSM_reg_3 ( .CK(PCICLK), .D(ITDSMNXT_3), .R(TRST_), .Q(ITDSM[3])
         );
    zivb U1033 ( .A(n2120), .Y(ITDSMNXT_7) );
    zivb U1034 ( .A(ITDSM[7]), .Y(n1846) );
    zbfb U1035 ( .A(n1993), .Y(n1769) );
    zbfb U1036 ( .A(DW9[8]), .Y(TRAN_CMD[29]) );
    zbfb U1037 ( .A(DW9[9]), .Y(TRAN_CMD[30]) );
    zbfb U1038 ( .A(DW9[10]), .Y(TRAN_CMD[31]) );
    zbfb U1039 ( .A(DW9[11]), .Y(TRAN_CMD[32]) );
    zbfb U1040 ( .A(DW9[0]), .Y(TRAN_CMD[33]) );
    zbfb U1041 ( .A(DW9[1]), .Y(TRAN_CMD[34]) );
    zbfb U1042 ( .A(DW9[2]), .Y(TRAN_CMD[35]) );
    zbfb U1043 ( .A(DW9[3]), .Y(TRAN_CMD[36]) );
    zbfb U1044 ( .A(DW9[4]), .Y(TRAN_CMD[37]) );
    zbfb U1045 ( .A(DW9[5]), .Y(TRAN_CMD[38]) );
    zbfb U1046 ( .A(DW9[6]), .Y(TRAN_CMD[39]) );
    zivb U1047 ( .A(n2203), .Y(TRAN_CMD[104]) );
    zbfb U1048 ( .A(IHCIADD[28]), .Y(IRXERR) );
    zdffqrb_ IRXERR_reg ( .CK(PCICLK), .D(IRXERR1209), .R(TRST_), .Q(IHCIADD
        [28]) );
    zbfb U1049 ( .A(BABBLE), .Y(IHCIADD[29]) );
    zivb U1050 ( .A(n1759), .Y(IHCIREQ) );
    zbfb U1051 ( .A(ITDSM[0]), .Y(ITDIDLE) );
    zdffsb ITDSM_reg_0 ( .CK(PCICLK), .D(PHASENXT_idle), .S(TRST_), .Q(ITDSM
        [0]), .QN(n1869) );
    zxo2b U1052 ( .A(add_487_carry_29), .B(CACHE_ADDR[26]), .Y(IHCIADR[31]) );
    zan2b U1053 ( .A(CACHE_ADDR[25]), .B(add_487_carry_28), .Y(
        add_487_carry_29) );
    zxo2b U1054 ( .A(CACHE_ADDR[25]), .B(add_487_carry_28), .Y(IHCIADR[30]) );
    zan2b U1055 ( .A(CACHE_ADDR[24]), .B(add_487_carry_27), .Y(
        add_487_carry_28) );
    zxo2b U1056 ( .A(CACHE_ADDR[24]), .B(add_487_carry_27), .Y(IHCIADR[29]) );
    zan2b U1057 ( .A(CACHE_ADDR[23]), .B(add_487_carry_26), .Y(
        add_487_carry_27) );
    zxo2b U1058 ( .A(CACHE_ADDR[23]), .B(add_487_carry_26), .Y(IHCIADR[28]) );
    zan2b U1059 ( .A(CACHE_ADDR[22]), .B(add_487_carry_25), .Y(
        add_487_carry_26) );
    zxo2b U1060 ( .A(CACHE_ADDR[22]), .B(add_487_carry_25), .Y(IHCIADR[27]) );
    zan2b U1061 ( .A(CACHE_ADDR[21]), .B(add_487_carry_24), .Y(
        add_487_carry_25) );
    zxo2b U1062 ( .A(CACHE_ADDR[21]), .B(add_487_carry_24), .Y(IHCIADR[26]) );
    zan2b U1063 ( .A(CACHE_ADDR[20]), .B(add_487_carry_23), .Y(
        add_487_carry_24) );
    zxo2b U1064 ( .A(CACHE_ADDR[20]), .B(add_487_carry_23), .Y(IHCIADR[25]) );
    zan2b U1065 ( .A(CACHE_ADDR[19]), .B(add_487_carry_22), .Y(
        add_487_carry_23) );
    zxo2b U1066 ( .A(CACHE_ADDR[19]), .B(add_487_carry_22), .Y(IHCIADR[24]) );
    zan2b U1067 ( .A(CACHE_ADDR[18]), .B(add_487_carry_21), .Y(
        add_487_carry_22) );
    zxo2b U1068 ( .A(CACHE_ADDR[18]), .B(add_487_carry_21), .Y(IHCIADR[23]) );
    zan2b U1069 ( .A(CACHE_ADDR[17]), .B(add_487_carry_20), .Y(
        add_487_carry_21) );
    zxo2b U1070 ( .A(CACHE_ADDR[17]), .B(add_487_carry_20), .Y(IHCIADR[22]) );
    zan2b U1071 ( .A(CACHE_ADDR[16]), .B(add_487_carry_19), .Y(
        add_487_carry_20) );
    zxo2b U1072 ( .A(CACHE_ADDR[16]), .B(add_487_carry_19), .Y(IHCIADR[21]) );
    zan2b U1073 ( .A(CACHE_ADDR[15]), .B(add_487_carry_18), .Y(
        add_487_carry_19) );
    zxo2b U1074 ( .A(CACHE_ADDR[15]), .B(add_487_carry_18), .Y(IHCIADR[20]) );
    zan2b U1075 ( .A(CACHE_ADDR[14]), .B(add_487_carry_17), .Y(
        add_487_carry_18) );
    zxo2b U1076 ( .A(CACHE_ADDR[14]), .B(add_487_carry_17), .Y(IHCIADR[19]) );
    zan2b U1077 ( .A(CACHE_ADDR[13]), .B(add_487_carry_16), .Y(
        add_487_carry_17) );
    zxo2b U1078 ( .A(CACHE_ADDR[13]), .B(add_487_carry_16), .Y(IHCIADR[18]) );
    zan2b U1079 ( .A(CACHE_ADDR[12]), .B(add_487_carry_15), .Y(
        add_487_carry_16) );
    zxo2b U1080 ( .A(CACHE_ADDR[12]), .B(add_487_carry_15), .Y(IHCIADR[17]) );
    zan2b U1081 ( .A(CACHE_ADDR[11]), .B(add_487_carry_14), .Y(
        add_487_carry_15) );
    zxo2b U1082 ( .A(CACHE_ADDR[11]), .B(add_487_carry_14), .Y(IHCIADR[16]) );
    zan2b U1083 ( .A(CACHE_ADDR[10]), .B(add_487_carry_13), .Y(
        add_487_carry_14) );
    zxo2b U1084 ( .A(CACHE_ADDR[10]), .B(add_487_carry_13), .Y(IHCIADR[15]) );
    zan2b U1085 ( .A(CACHE_ADDR[9]), .B(add_487_carry_12), .Y(add_487_carry_13
        ) );
    zxo2b U1086 ( .A(CACHE_ADDR[9]), .B(add_487_carry_12), .Y(IHCIADR[14]) );
    zan2b U1087 ( .A(CACHE_ADDR[8]), .B(add_487_carry_11), .Y(add_487_carry_12
        ) );
    zxo2b U1088 ( .A(CACHE_ADDR[8]), .B(add_487_carry_11), .Y(IHCIADR[13]) );
    zan2b U1089 ( .A(CACHE_ADDR[7]), .B(add_487_carry_10), .Y(add_487_carry_11
        ) );
    zxo2b U1090 ( .A(CACHE_ADDR[7]), .B(add_487_carry_10), .Y(IHCIADR[12]) );
    zan2b U1091 ( .A(CACHE_ADDR[6]), .B(add_487_carry_9), .Y(add_487_carry_10)
         );
    zxo2b U1092 ( .A(CACHE_ADDR[6]), .B(add_487_carry_9), .Y(IHCIADR[11]) );
    zan2b U1093 ( .A(CACHE_ADDR[5]), .B(add_487_carry_8), .Y(add_487_carry_9)
         );
    zxo2b U1094 ( .A(CACHE_ADDR[5]), .B(add_487_carry_8), .Y(IHCIADR[10]) );
    zan2b U1095 ( .A(CACHE_ADDR[4]), .B(add_487_carry_7), .Y(add_487_carry_8)
         );
    zxo2b U1096 ( .A(CACHE_ADDR[4]), .B(add_487_carry_7), .Y(IHCIADR[9]) );
    zan2b U1097 ( .A(CACHE_ADDR[3]), .B(add_487_carry_6), .Y(add_487_carry_7)
         );
    zxo2b U1098 ( .A(CACHE_ADDR[3]), .B(add_487_carry_6), .Y(IHCIADR[8]) );
    zan2b U1099 ( .A(CACHE_ADDR[2]), .B(add_487_carry_5), .Y(add_487_carry_6)
         );
    zxo2b U1100 ( .A(CACHE_ADDR[2]), .B(add_487_carry_5), .Y(IHCIADR[7]) );
    zan2b U1101 ( .A(CACHE_ADDR[1]), .B(add_487_carry_4), .Y(add_487_carry_5)
         );
    zxo2b U1102 ( .A(CACHE_ADDR[1]), .B(add_487_carry_4), .Y(IHCIADR[6]) );
    zan2b U1103 ( .A(CACHE_ADDR[0]), .B(add_487_carry_3), .Y(add_487_carry_4)
         );
    zxo2b U1104 ( .A(CACHE_ADDR[0]), .B(add_487_carry_3), .Y(IHCIADR[5]) );
    zan2b U1105 ( .A(FRNUM[2]), .B(add_487_carry_2), .Y(add_487_carry_3) );
    zxo2b U1106 ( .A(FRNUM[2]), .B(add_487_carry_2), .Y(IHCIADR[4]) );
    zan2b U1107 ( .A(FRNUM[1]), .B(FRNUM[0]), .Y(add_487_carry_2) );
    zxo2b U1108 ( .A(FRNUM[1]), .B(FRNUM[0]), .Y(IHCIADR[3]) );
    zxn2b U1109 ( .A(sub_328_carry_11), .B(TRANSLEN_11), .Y(TRANSLEN795_11) );
    zor2b U1110 ( .A(TRANSLEN_0), .B(sub_328_B_not_0), .Y(sub_328_carry_1) );
    zxn2b U1111 ( .A(TRANSLEN_0), .B(sub_328_B_not_0), .Y(TRANSLEN795_0) );
    zxo2b U1112 ( .A(add_353_carry_11), .B(TR_LEN_11), .Y(TR_LEN913_11) );
    zan2b U1113 ( .A(TR_LEN_0), .B(ACTLEN[0]), .Y(add_353_carry_1) );
    zxo2b U1114 ( .A(TR_LEN_0), .B(ACTLEN[0]), .Y(TR_LEN913_0) );
    zxo2b U1115 ( .A(r211_carry_12), .B(TRANSOFFSET_12), .Y(TRANSOFFSET1141_12
        ) );
    zan2b U1116 ( .A(TRAN_CMD[83]), .B(r211_carry_11), .Y(r211_carry_12) );
    zxo2b U1117 ( .A(TRAN_CMD[83]), .B(r211_carry_11), .Y(TRANSOFFSET1141_11)
         );
    zan2b U1118 ( .A(_cell_414_U49_Z_0), .B(TRAN_CMD[72]), .Y(r211_carry_1) );
    zxo2b U1119 ( .A(_cell_414_U49_Z_0), .B(TRAN_CMD[72]), .Y(
        TRANSOFFSET1141_0) );
    zdffrb ITDSM_reg_11 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(ITDSM[11]) );
    zdffrb ITDSM_reg_10 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(ITDSM[10]) );
    zdffrb ITDSM_reg_12 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(ITDSM[12]) );
    zdffrb ITDSM_reg_13 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(ITDSM[13]) );
    znd2d U1124 ( .A(n1839), .B(n1758), .Y(LENGTMAX_PRE) );
    zfa1b sub_328_U2_6 ( .A(TRANSLEN_6), .B(sub_328_B_not_6), .CI(
        sub_328_carry_6), .CO(sub_328_carry_7), .S(TRANSLEN795_6) );
    zfa1b sub_328_U2_8 ( .A(TRANSLEN_8), .B(sub_328_B_not_8), .CI(
        sub_328_carry_8), .CO(sub_328_carry_9), .S(TRANSLEN795_8) );
    zfa1b sub_328_U2_10 ( .A(TRANSLEN_10), .B(sub_328_B_not_10), .CI(
        sub_328_carry_10), .CO(sub_328_carry_11), .S(TRANSLEN795_10) );
    zfa1b sub_328_U2_9 ( .A(TRANSLEN_9), .B(sub_328_B_not_9), .CI(
        sub_328_carry_9), .CO(sub_328_carry_10), .S(TRANSLEN795_9) );
    zfa1b sub_328_U2_1 ( .A(TRANSLEN_1), .B(sub_328_B_not_1), .CI(
        sub_328_carry_1), .CO(sub_328_carry_2), .S(TRANSLEN795_1) );
    zfa1b sub_328_U2_7 ( .A(TRANSLEN_7), .B(sub_328_B_not_7), .CI(
        sub_328_carry_7), .CO(sub_328_carry_8), .S(TRANSLEN795_7) );
    zfa1b sub_328_U2_5 ( .A(TRANSLEN_5), .B(sub_328_B_not_5), .CI(
        sub_328_carry_5), .CO(sub_328_carry_6), .S(TRANSLEN795_5) );
    zfa1b sub_328_U2_3 ( .A(TRANSLEN_3), .B(sub_328_B_not_3), .CI(
        sub_328_carry_3), .CO(sub_328_carry_4), .S(TRANSLEN795_3) );
    zfa1b sub_328_U2_2 ( .A(TRANSLEN_2), .B(sub_328_B_not_2), .CI(
        sub_328_carry_2), .CO(sub_328_carry_3), .S(TRANSLEN795_2) );
    zfa1b sub_328_U2_4 ( .A(TRANSLEN_4), .B(sub_328_B_not_4), .CI(
        sub_328_carry_4), .CO(sub_328_carry_5), .S(TRANSLEN795_4) );
    zfa1b add_353_U1_5 ( .A(ACTLEN[5]), .B(TR_LEN_5), .CI(add_353_carry_5), 
        .CO(add_353_carry_6), .S(TR_LEN913_5) );
    zfa1b add_353_U1_4 ( .A(ACTLEN[4]), .B(TR_LEN_4), .CI(add_353_carry_4), 
        .CO(add_353_carry_5), .S(TR_LEN913_4) );
    zfa1b add_353_U1_3 ( .A(ACTLEN[3]), .B(TR_LEN_3), .CI(add_353_carry_3), 
        .CO(add_353_carry_4), .S(TR_LEN913_3) );
    zfa1b add_353_U1_10 ( .A(ACTLEN[10]), .B(TR_LEN_10), .CI(add_353_carry_10), 
        .CO(add_353_carry_11), .S(TR_LEN913_10) );
    zfa1b add_353_U1_9 ( .A(ACTLEN[9]), .B(TR_LEN_9), .CI(add_353_carry_9), 
        .CO(add_353_carry_10), .S(TR_LEN913_9) );
    zfa1b add_353_U1_2 ( .A(ACTLEN[2]), .B(TR_LEN_2), .CI(add_353_carry_2), 
        .CO(add_353_carry_3), .S(TR_LEN913_2) );
    zfa1b add_353_U1_7 ( .A(ACTLEN[7]), .B(TR_LEN_7), .CI(add_353_carry_7), 
        .CO(add_353_carry_8), .S(TR_LEN913_7) );
    zfa1b add_353_U1_8 ( .A(ACTLEN[8]), .B(TR_LEN_8), .CI(add_353_carry_8), 
        .CO(add_353_carry_9), .S(TR_LEN913_8) );
    zfa1b add_353_U1_6 ( .A(ACTLEN[6]), .B(TR_LEN_6), .CI(add_353_carry_6), 
        .CO(add_353_carry_7), .S(TR_LEN913_6) );
    zfa1b add_353_U1_1 ( .A(ACTLEN[1]), .B(TR_LEN_1), .CI(add_353_carry_1), 
        .CO(add_353_carry_2), .S(TR_LEN913_1) );
    zfa1b r211_U1_5 ( .A(TRAN_CMD[77]), .B(_cell_414_U49_Z_5), .CI(
        r211_carry_5), .CO(r211_carry_6), .S(TRANSOFFSET1141_5) );
    zfa1b r211_U1_4 ( .A(TRAN_CMD[76]), .B(_cell_414_U49_Z_4), .CI(
        r211_carry_4), .CO(r211_carry_5), .S(TRANSOFFSET1141_4) );
    zfa1b r211_U1_3 ( .A(TRAN_CMD[75]), .B(_cell_414_U49_Z_3), .CI(
        r211_carry_3), .CO(r211_carry_4), .S(TRANSOFFSET1141_3) );
    zfa1b r211_U1_10 ( .A(TRAN_CMD[82]), .B(_cell_414_U49_Z_10), .CI(
        r211_carry_10), .CO(r211_carry_11), .S(TRANSOFFSET1141_10) );
    zfa1b r211_U1_9 ( .A(TRAN_CMD[81]), .B(_cell_414_U49_Z_9), .CI(
        r211_carry_9), .CO(r211_carry_10), .S(TRANSOFFSET1141_9) );
    zfa1b r211_U1_2 ( .A(TRAN_CMD[74]), .B(_cell_414_U49_Z_2), .CI(
        r211_carry_2), .CO(r211_carry_3), .S(TRANSOFFSET1141_2) );
    zfa1b r211_U1_7 ( .A(TRAN_CMD[79]), .B(_cell_414_U49_Z_7), .CI(
        r211_carry_7), .CO(r211_carry_8), .S(TRANSOFFSET1141_7) );
    zfa1b r211_U1_8 ( .A(TRAN_CMD[80]), .B(_cell_414_U49_Z_8), .CI(
        r211_carry_8), .CO(r211_carry_9), .S(TRANSOFFSET1141_8) );
    zfa1b r211_U1_6 ( .A(TRAN_CMD[78]), .B(_cell_414_U49_Z_6), .CI(
        r211_carry_6), .CO(r211_carry_7), .S(TRANSOFFSET1141_6) );
    zfa1b r211_U1_1 ( .A(TRAN_CMD[73]), .B(_cell_414_U49_Z_1), .CI(
        r211_carry_1), .CO(r211_carry_2), .S(TRANSOFFSET1141_1) );
    zao211b U1125 ( .A(n1737), .B(n1843), .C(n1844), .D(n1845), .Y(
        PHASENXT_idle) );
    zoa21d U1126 ( .A(ICMDSTART_EOT), .B(ICMDSTART), .C(n1857), .Y(
        ICMDSTART_EOT1246) );
    zao211b U1127 ( .A(n1862), .B(n1863), .C(ITDSM[6]), .D(n1864), .Y(IEOT1283
        ) );
    zoa21d U1128 ( .A(PG_INC), .B(TRANSOFFSET_12), .C(n1870), .Y(PG_INC472) );
    zao222b U1129 ( .A(TRANSLEN795_11), .B(n1873), .C(n1874), .D(n1875), .E(
        TRANSLEN_11), .F(n1876), .Y(TRANSLEN813_11) );
    zao222b U1130 ( .A(TRANSLEN795_10), .B(n1873), .C(LDPARM), .D(n1877), .E(
        TRANSLEN_10), .F(n1876), .Y(TRANSLEN813_10) );
    zao222b U1131 ( .A(n1873), .B(TRANSLEN795_9), .C(n1874), .D(n1878), .E(
        TRANSLEN_9), .F(n1876), .Y(TRANSLEN813_9) );
    zao222b U1132 ( .A(TRANSLEN795_8), .B(n1873), .C(LDPARM), .D(n1879), .E(
        TRANSLEN_8), .F(n1876), .Y(TRANSLEN813_8) );
    zao222b U1133 ( .A(TRANSLEN795_7), .B(n1873), .C(n1874), .D(n1880), .E(
        TRANSLEN_7), .F(n1876), .Y(TRANSLEN813_7) );
    zao222b U1134 ( .A(TRANSLEN795_6), .B(n1873), .C(LDPARM), .D(n1881), .E(
        TRANSLEN_6), .F(n1876), .Y(TRANSLEN813_6) );
    zao222b U1135 ( .A(TRANSLEN795_5), .B(n1873), .C(n1874), .D(n1882), .E(
        TRANSLEN_5), .F(n1876), .Y(TRANSLEN813_5) );
    zao222b U1136 ( .A(TRANSLEN795_4), .B(n1873), .C(LDPARM), .D(n1883), .E(
        TRANSLEN_4), .F(n1876), .Y(TRANSLEN813_4) );
    zao222b U1137 ( .A(TRANSLEN795_3), .B(n1873), .C(n1874), .D(n1884), .E(
        TRANSLEN_3), .F(n1876), .Y(TRANSLEN813_3) );
    zao222b U1138 ( .A(TRANSLEN795_2), .B(n1873), .C(LDPARM), .D(n1885), .E(
        TRANSLEN_2), .F(n1876), .Y(TRANSLEN813_2) );
    zao222b U1139 ( .A(TRANSLEN795_1), .B(n1873), .C(n1874), .D(n1886), .E(
        TRANSLEN_1), .F(n1876), .Y(TRANSLEN813_1) );
    zao222b U1140 ( .A(TRANSLEN795_0), .B(n1873), .C(LDPARM), .D(n1887), .E(
        TRANSLEN_0), .F(n1876), .Y(TRANSLEN813_0) );
    zao211b U1141 ( .A(n1016), .B(n1891), .C(n1892), .D(n1893), .Y(MULT612_1)
         );
    zao222b U1142 ( .A(n1874), .B(DW11[0]), .C(n1894), .D(NXTISSTSWB), .E(
        MULT_0), .F(n1891), .Y(MULT612_0) );
    zao222b U1143 ( .A(LDPARM), .B(IHCIADD[11]), .C(TRAN_CMD[83]), .D(n1891), 
        .E(TRANSOFFSET1141_11), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_11) );
    zao222b U1144 ( .A(n1874), .B(IHCIADD[10]), .C(TRAN_CMD[82]), .D(n1891), 
        .E(TRANSOFFSET1141_10), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_10) );
    zao222b U1145 ( .A(LDPARM), .B(IHCIADD[9]), .C(TRAN_CMD[81]), .D(n1891), 
        .E(TRANSOFFSET1141_9), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_9) );
    zao222b U1146 ( .A(n1874), .B(IHCIADD[8]), .C(TRAN_CMD[80]), .D(n1891), 
        .E(TRANSOFFSET1141_8), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_8) );
    zao222b U1147 ( .A(LDPARM), .B(IHCIADD[7]), .C(TRAN_CMD[79]), .D(n1891), 
        .E(TRANSOFFSET1141_7), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_7) );
    zao222b U1148 ( .A(n1874), .B(IHCIADD[6]), .C(TRAN_CMD[78]), .D(n1891), 
        .E(TRANSOFFSET1141_6), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_6) );
    zao222b U1149 ( .A(LDPARM), .B(IHCIADD[5]), .C(TRAN_CMD[77]), .D(n1891), 
        .E(TRANSOFFSET1141_5), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_5) );
    zao222b U1150 ( .A(n1874), .B(IHCIADD[4]), .C(TRAN_CMD[76]), .D(n1891), 
        .E(TRANSOFFSET1141_4), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_4) );
    zao222b U1151 ( .A(LDPARM), .B(IHCIADD[3]), .C(TRAN_CMD[75]), .D(n1891), 
        .E(TRANSOFFSET1141_3), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_3) );
    zao222b U1152 ( .A(n1874), .B(IHCIADD[2]), .C(TRAN_CMD[74]), .D(n1891), 
        .E(TRANSOFFSET1141_2), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_2) );
    zao222b U1153 ( .A(LDPARM), .B(IHCIADD[1]), .C(TRAN_CMD[73]), .D(n1891), 
        .E(TRANSOFFSET1141_1), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_1) );
    zao222b U1154 ( .A(n1874), .B(IHCIADD[0]), .C(TRAN_CMD[72]), .D(n1891), 
        .E(TRANSOFFSET1141_0), .F(NXTISSTSWB), .Y(TRANSOFFSET1140_0) );
    zao211b U1155 ( .A(ITDSM[9]), .B(n1921), .C(GEN_PERR), .D(n1922), .Y(
        ITDERRINT_T1513) );
    zan4b U1156 ( .A(n1869), .B(n1888), .C(n1923), .D(n1924), .Y(IRXERR1209)
         );
    zor3b U1157 ( .A(n1933), .B(n1934), .C(n1935), .Y(TRAN_CMD[103]) );
    zor3b U1158 ( .A(n1936), .B(n1937), .C(n1938), .Y(TRAN_CMD[102]) );
    zor3b U1159 ( .A(n1939), .B(n1940), .C(n1941), .Y(TRAN_CMD[101]) );
    zor3b U1160 ( .A(n1942), .B(n1943), .C(n1944), .Y(TRAN_CMD[100]) );
    zor3b U1161 ( .A(n1945), .B(n1946), .C(n1947), .Y(TRAN_CMD[99]) );
    zor3b U1162 ( .A(n1948), .B(n1949), .C(n1950), .Y(TRAN_CMD[98]) );
    zor3b U1163 ( .A(n1951), .B(n1952), .C(n1953), .Y(TRAN_CMD[97]) );
    zor3b U1164 ( .A(n1954), .B(n1955), .C(n1956), .Y(TRAN_CMD[96]) );
    zor3b U1165 ( .A(n1957), .B(n1958), .C(n1959), .Y(TRAN_CMD[95]) );
    zor3b U1166 ( .A(n1960), .B(n1961), .C(n1962), .Y(TRAN_CMD[94]) );
    zor3b U1167 ( .A(n1963), .B(n1964), .C(n1965), .Y(TRAN_CMD[93]) );
    zor3b U1168 ( .A(n1966), .B(n1967), .C(n1968), .Y(TRAN_CMD[92]) );
    zor3b U1169 ( .A(n1969), .B(n1970), .C(n1971), .Y(TRAN_CMD[91]) );
    zor3b U1170 ( .A(n1972), .B(n1973), .C(n1974), .Y(TRAN_CMD[90]) );
    zor3b U1171 ( .A(n1975), .B(n1976), .C(n1977), .Y(TRAN_CMD[89]) );
    zor3b U1172 ( .A(n1978), .B(n1979), .C(n1980), .Y(TRAN_CMD[88]) );
    zor3b U1173 ( .A(n1981), .B(n1982), .C(n1983), .Y(TRAN_CMD[87]) );
    zor3b U1174 ( .A(n1984), .B(n1985), .C(n1986), .Y(TRAN_CMD[86]) );
    zor3b U1175 ( .A(n1987), .B(n1988), .C(n1989), .Y(TRAN_CMD[85]) );
    zor3b U1176 ( .A(n1990), .B(n1991), .C(n1992), .Y(TRAN_CMD[84]) );
    zao211b U1177 ( .A(DW15[12]), .B(n1993), .C(n1994), .D(n1995), .Y(TRAN_CMD
        [52]) );
    zao211b U1178 ( .A(DW15[13]), .B(n1993), .C(n1996), .D(n1997), .Y(TRAN_CMD
        [53]) );
    zao211b U1179 ( .A(DW15[14]), .B(n1993), .C(n1998), .D(n1999), .Y(TRAN_CMD
        [54]) );
    zao211b U1180 ( .A(DW15[15]), .B(n1769), .C(n2000), .D(n2001), .Y(TRAN_CMD
        [55]) );
    zao211b U1181 ( .A(DW15[16]), .B(n1993), .C(n2002), .D(n2003), .Y(TRAN_CMD
        [56]) );
    zao211b U1182 ( .A(DW15[17]), .B(n1993), .C(n2004), .D(n2005), .Y(TRAN_CMD
        [57]) );
    zao211b U1183 ( .A(DW15[18]), .B(n1993), .C(n2006), .D(n2007), .Y(TRAN_CMD
        [58]) );
    zao211b U1184 ( .A(DW15[19]), .B(n1993), .C(n2008), .D(n2009), .Y(TRAN_CMD
        [59]) );
    zao211b U1185 ( .A(DW15[20]), .B(n1993), .C(n2010), .D(n2011), .Y(TRAN_CMD
        [60]) );
    zao211b U1186 ( .A(DW15[21]), .B(n1993), .C(n2012), .D(n2013), .Y(TRAN_CMD
        [61]) );
    zao211b U1187 ( .A(DW15[22]), .B(n1769), .C(n2014), .D(n2015), .Y(TRAN_CMD
        [62]) );
    zao211b U1188 ( .A(DW15[23]), .B(n1769), .C(n2016), .D(n2017), .Y(TRAN_CMD
        [63]) );
    zao211b U1189 ( .A(DW15[24]), .B(n1993), .C(n2018), .D(n2019), .Y(TRAN_CMD
        [64]) );
    zao211b U1190 ( .A(DW15[25]), .B(n1993), .C(n2020), .D(n2021), .Y(TRAN_CMD
        [65]) );
    zao211b U1191 ( .A(DW15[26]), .B(n1993), .C(n2022), .D(n2023), .Y(TRAN_CMD
        [66]) );
    zao211b U1192 ( .A(DW15[27]), .B(n1993), .C(n2024), .D(n2025), .Y(TRAN_CMD
        [67]) );
    zao211b U1193 ( .A(DW15[28]), .B(n1769), .C(n2026), .D(n2027), .Y(TRAN_CMD
        [68]) );
    zao211b U1194 ( .A(DW15[29]), .B(n1769), .C(n2028), .D(n2029), .Y(TRAN_CMD
        [69]) );
    zao211b U1195 ( .A(DW15[30]), .B(n1993), .C(n2030), .D(n2031), .Y(TRAN_CMD
        [70]) );
    zao211b U1196 ( .A(DW15[31]), .B(n1993), .C(n2032), .D(n2033), .Y(TRAN_CMD
        [71]) );
    zoa21d U1197 ( .A(RXDATA0), .B(SPD), .C(TRAN_CMD[104]), .Y(n2039) );
    zoa21d U1198 ( .A(DW11[1]), .B(n1925), .C(TRAN_CMD[8]), .Y(n2045) );
    zcx8d U1199 ( .A(n2045), .B(n2048), .C(n2041), .D(n2047), .E(n2201), .Y(
        n2046) );
    zoa21d U1200 ( .A(IHCIADD[28]), .B(n2053), .C(n1858), .Y(n2052) );
    zoa21d U1201 ( .A(RXDATA2), .B(RXDATA0), .C(n2201), .Y(n2058) );
    zan4b U1202 ( .A(n1735), .B(MULT650_1), .C(n2060), .D(NXTISSTSWB), .Y(
        n1892) );
    zoa21d U1203 ( .A(n2066), .B(n2067), .C(ITDSM[9]), .Y(n2065) );
    zor4b U1204 ( .A(ITDSM[11]), .B(ITDSM[10]), .C(ITDSM[13]), .D(ITDSM[12]), 
        .Y(n2068) );
    zor4b U1205 ( .A(ITDSM[9]), .B(ITDSM[7]), .C(ITDSM[5]), .D(n2068), .Y(
        n2069) );
    zor3b U1206 ( .A(ITDSM[6]), .B(ITDSM[8]), .C(n2069), .Y(n2070) );
    zor3b U1207 ( .A(IHCIADR[2]), .B(n2073), .C(n2074), .Y(n2075) );
    zor3b U1208 ( .A(FRNUM[0]), .B(n2073), .C(n2074), .Y(n2076) );
    zor3b U1209 ( .A(FRNUM[1]), .B(IHCIADR[2]), .C(n2074), .Y(n2077) );
    zor3b U1210 ( .A(FRNUM[1]), .B(FRNUM[0]), .C(n2074), .Y(n2078) );
    zor3b U1211 ( .A(FRNUM[2]), .B(IHCIADR[2]), .C(n2073), .Y(n2079) );
    zor3b U1212 ( .A(FRNUM[2]), .B(FRNUM[0]), .C(n2073), .Y(n2080) );
    zor3b U1213 ( .A(FRNUM[2]), .B(FRNUM[1]), .C(IHCIADR[2]), .Y(n2081) );
    zor3b U1214 ( .A(FRNUM[2]), .B(FRNUM[1]), .C(FRNUM[0]), .Y(n2082) );
    zor4b U1215 ( .A(n2040), .B(n1870), .C(RECOVERYMODE), .D(n2083), .Y(n1843)
         );
    zor3b U1216 ( .A(ITDSM[3]), .B(n2084), .C(n1863), .Y(n2056) );
    zor4b U1217 ( .A(n1862), .B(n2086), .C(n2088), .D(n2039), .Y(n2087) );
    zor4b U1218 ( .A(ITDSM[0]), .B(n1863), .C(n2038), .D(n2071), .Y(n2089) );
    zor3b U1219 ( .A(PG_1), .B(n2109), .C(n2106), .Y(n2110) );
    zor3b U1220 ( .A(PG_1), .B(PG_0), .C(n2106), .Y(n2111) );
    zor3b U1221 ( .A(n2109), .B(n2107), .C(PG_2), .Y(n2112) );
    zor3b U1222 ( .A(n2107), .B(PG_0), .C(PG_2), .Y(n2113) );
    zor3b U1223 ( .A(PG_1), .B(n2109), .C(PG_2), .Y(n2114) );
    zor3b U1224 ( .A(PG_1), .B(PG_0), .C(PG_2), .Y(n2115) );
    zor3b U1225 ( .A(n2069), .B(n2092), .C(n2066), .Y(n2050) );
    zor3b U1226 ( .A(ITDSM[6]), .B(n2068), .C(n2066), .Y(n2119) );
    zor4b U1227 ( .A(ITDSM[9]), .B(ITDSM[5]), .C(n1846), .D(n2119), .Y(n2051)
         );
    zor3b U1228 ( .A(IHCIADD[28]), .B(n1765), .C(n2053), .Y(n2123) );
    zor3b U1229 ( .A(n1857), .B(n2089), .C(GEN_PERR), .Y(n2130) );
    zaoi2x4d U1230 ( .A(n2204), .B(DW8[31]), .C(n2175), .D(DW7[31]), .E(n2176), 
        .F(DW6[31]), .G(n2177), .H(DW5[31]), .Y(n1866) );
    zao222b U1231 ( .A(n2186), .B(DW10[27]), .C(n2213), .D(DW11[27]), .E(n2214
        ), .F(DW9[27]), .Y(n1946) );
    zao222b U1232 ( .A(DW10[26]), .B(n2212), .C(DW11[26]), .D(n2213), .E(DW9
        [26]), .F(n2214), .Y(n1949) );
    zao222b U1233 ( .A(DW10[25]), .B(n2186), .C(DW11[25]), .D(n2187), .E(DW9
        [25]), .F(n2188), .Y(n1952) );
    zao222b U1234 ( .A(DW10[24]), .B(n2212), .C(DW11[24]), .D(n2213), .E(DW9
        [24]), .F(n2214), .Y(n1955) );
    zao222b U1235 ( .A(DW10[23]), .B(n2186), .C(DW11[23]), .D(n2187), .E(DW9
        [23]), .F(n2188), .Y(n1958) );
    zao222b U1236 ( .A(DW10[22]), .B(n2212), .C(DW11[22]), .D(n2213), .E(DW9
        [22]), .F(n2214), .Y(n1961) );
    zao222b U1237 ( .A(DW10[21]), .B(n2186), .C(DW11[21]), .D(n2187), .E(DW9
        [21]), .F(n2188), .Y(n1964) );
    zao222b U1238 ( .A(DW10[20]), .B(n2212), .C(DW11[20]), .D(n2213), .E(DW9
        [20]), .F(n2214), .Y(n1967) );
    zao222b U1239 ( .A(DW10[19]), .B(n2186), .C(DW11[19]), .D(n2187), .E(DW9
        [19]), .F(n2188), .Y(n1970) );
    zao222b U1240 ( .A(DW10[18]), .B(n2212), .C(DW11[18]), .D(n2213), .E(DW9
        [18]), .F(n2214), .Y(n1973) );
    zao222b U1241 ( .A(DW10[17]), .B(n2186), .C(DW11[17]), .D(n2187), .E(DW9
        [17]), .F(n2188), .Y(n1976) );
    zao222b U1242 ( .A(DW10[16]), .B(n2186), .C(DW11[16]), .D(n2213), .E(DW9
        [16]), .F(n2214), .Y(n1979) );
    zao222b U1243 ( .A(DW10[15]), .B(n2212), .C(DW11[15]), .D(n2187), .E(DW9
        [15]), .F(n2188), .Y(n1982) );
    zao222b U1244 ( .A(DW10[14]), .B(n2212), .C(DW11[14]), .D(n2213), .E(DW9
        [14]), .F(n2214), .Y(n1985) );
    zao222b U1245 ( .A(DW10[13]), .B(n2186), .C(DW11[13]), .D(n2187), .E(DW9
        [13]), .F(n2188), .Y(n1988) );
    zao222b U1246 ( .A(DW10[12]), .B(n2212), .C(DW11[12]), .D(n2213), .E(DW9
        [12]), .F(n2214), .Y(n1991) );
    zao222b U1247 ( .A(DW11[31]), .B(n2186), .C(DW12[31]), .D(n2187), .E(DW10
        [31]), .F(n2188), .Y(n2032) );
    zao222b U1248 ( .A(DW11[30]), .B(n2212), .C(DW12[30]), .D(n2213), .E(DW10
        [30]), .F(n2188), .Y(n2030) );
    zao222b U1249 ( .A(DW11[29]), .B(n2186), .C(DW12[29]), .D(n2187), .E(DW10
        [29]), .F(n2214), .Y(n2028) );
    zao222b U1250 ( .A(DW11[28]), .B(n2212), .C(DW12[28]), .D(n2213), .E(DW10
        [28]), .F(n2188), .Y(n2026) );
    zao222b U1251 ( .A(n2212), .B(DW11[27]), .C(n2187), .D(DW12[27]), .E(n2188
        ), .F(DW10[27]), .Y(n2024) );
    zao222b U1252 ( .A(DW11[26]), .B(n2186), .C(DW12[26]), .D(n2187), .E(DW10
        [26]), .F(n2214), .Y(n2022) );
    zao222b U1253 ( .A(DW11[25]), .B(n2212), .C(DW12[25]), .D(n2213), .E(DW10
        [25]), .F(n2214), .Y(n2020) );
    zao222b U1254 ( .A(DW11[24]), .B(n2186), .C(DW12[24]), .D(n2187), .E(DW10
        [24]), .F(n2188), .Y(n2018) );
    zao222b U1255 ( .A(DW11[23]), .B(n2212), .C(DW12[23]), .D(n2213), .E(DW10
        [23]), .F(n2214), .Y(n2016) );
    zao222b U1256 ( .A(DW11[22]), .B(n2186), .C(DW12[22]), .D(n2187), .E(DW10
        [22]), .F(n2188), .Y(n2014) );
    zao222b U1257 ( .A(DW11[21]), .B(n2212), .C(DW12[21]), .D(n2213), .E(DW10
        [21]), .F(n2214), .Y(n2012) );
    zao222b U1258 ( .A(DW11[20]), .B(n2186), .C(DW12[20]), .D(n2187), .E(DW10
        [20]), .F(n2188), .Y(n2010) );
    zao222b U1259 ( .A(DW11[19]), .B(n2212), .C(DW12[19]), .D(n2213), .E(DW10
        [19]), .F(n2214), .Y(n2008) );
    zao222b U1260 ( .A(DW11[18]), .B(n2186), .C(DW12[18]), .D(n2187), .E(DW10
        [18]), .F(n2188), .Y(n2006) );
    zao222b U1261 ( .A(DW11[17]), .B(n2212), .C(DW12[17]), .D(n2213), .E(DW10
        [17]), .F(n2214), .Y(n2004) );
    zao222b U1262 ( .A(DW11[16]), .B(n2186), .C(DW12[16]), .D(n2187), .E(DW10
        [16]), .F(n2188), .Y(n2002) );
    zao222b U1263 ( .A(DW11[15]), .B(n2212), .C(DW12[15]), .D(n2213), .E(DW10
        [15]), .F(n2188), .Y(n2000) );
    zao222b U1264 ( .A(DW11[14]), .B(n2186), .C(DW12[14]), .D(n2187), .E(DW10
        [14]), .F(n2214), .Y(n1998) );
    zao222b U1265 ( .A(DW11[13]), .B(n2212), .C(DW12[13]), .D(n2213), .E(DW10
        [13]), .F(n2214), .Y(n1996) );
    zao222b U1266 ( .A(DW11[12]), .B(n2186), .C(DW12[12]), .D(n2187), .E(DW10
        [12]), .F(n2188), .Y(n1994) );
    zao222b U1267 ( .A(DW10[31]), .B(n2212), .C(DW11[31]), .D(n2213), .E(DW9
        [31]), .F(n2214), .Y(n1934) );
    zao222b U1268 ( .A(DW10[30]), .B(n2186), .C(DW11[30]), .D(n2187), .E(DW9
        [30]), .F(n2188), .Y(n1937) );
    zao222b U1269 ( .A(DW10[29]), .B(n2186), .C(DW11[29]), .D(n2213), .E(DW9
        [29]), .F(n2188), .Y(n1940) );
    zao222b U1270 ( .A(DW10[28]), .B(n2212), .C(DW11[28]), .D(n2187), .E(DW9
        [28]), .F(n2214), .Y(n1943) );
    zao211b U1271 ( .A(ITDSM[7]), .B(n2126), .C(GEN_PERR), .D(n2189), .Y(n1844
        ) );
    zor4b U1272 ( .A(n2068), .B(n2134), .C(n2064), .D(n2065), .Y(n1845) );
    zor4b U1273 ( .A(PIDERR), .B(CRCERR), .C(TMOUT), .D(n2062), .Y(n2191) );
    zor6b U1274 ( .A(TRAN_CMD[47]), .B(TRAN_CMD[46]), .C(TRAN_CMD[45]), .D(
        TRAN_CMD[50]), .E(TRAN_CMD[49]), .F(TRAN_CMD[48]), .Y(n1853) );
    zor3b U1275 ( .A(ITDSM[4]), .B(ITDSM[5]), .C(n2063), .Y(n1860) );
    zao222b U1276 ( .A(n1742), .B(n2196), .C(n2194), .D(n1857), .E(n1737), .F(
        n2197), .Y(n2091) );
    zao21d U1277 ( .A(PG_0), .B(PG_2), .C(n2183), .Y(n1993) );
    zao222b U1278 ( .A(FEMPTY), .B(n2195), .C(n2198), .D(n1862), .E(n1739), 
        .F(n1890), .Y(n2122) );
    zor2d U1279 ( .A(n2052), .B(n1891), .Y(n1876) );
    zor3b U1280 ( .A(PARSEITDEND), .B(n1870), .C(n1856), .Y(n1859) );
    zao211b U1281 ( .A(n2200), .B(n2060), .C(n2191), .D(n2192), .Y(n2193) );
    zor3b U1282 ( .A(n2041), .B(n2116), .C(TRAN_CMD[8]), .Y(n2044) );
    zor3b U1283 ( .A(ITDSM[9]), .B(ITDSM[8]), .C(n2054), .Y(n2136) );
endmodule


module SITDCTL ( SITD_PARSE_GO, PARSESITDEND, SITDPARSING, SITDIDLE, FRNUM, 
    DW0, DW1, DW2, DW3, DW4, DW5, DW6, DW7, DW8, DW9, DW10, DW11, DW12, DW13, 
    GEN_PERR, PCIEND, DWCNT, CACHEPHASE, UP_DW3, UP_DW4, UP_DW5, UP_LDW3, 
    UP_LDW4, UP_LDW5, SIHCIREQ, SIDWNUM, SIDWOFFSET, SIHCIADR, SIHCIADD, 
    SIHCIMWR, SITDSM, TRAN_CMD, SITD_ACT, SIBUI_GO, CACHE_ADDR, CACHE_INVALID, 
    CRCERR, ACTLEN, BABBLE, PIDERR, TMOUT, RXDATA0, RXDATA1, RXMDATA, RXNYET, 
    RXPIDERR, EHCI_MAC_EOT, FEMPTY, TDMAEND, SIRXERR, SICMDSTART_REQ, 
    SICMDSTART, SIEOT, HCI_PRESOF, LTINT_PCLK, USBINT_EN, ERRINT_EN, USBINT, 
    ERRINT, SITDIOCINT_S, SITDERRINT_S, SITDIOCINT, RECOVERYMODE, PCICLK, 
    EHCIFLOW_PCLK, TRST_ );
input  [13:0] FRNUM;
input  [31:0] DW0;
output [31:0] SIHCIADD;
input  [31:0] DW7;
input  [31:0] DW9;
output [31:0] SIHCIADR;
input  [26:0] CACHE_ADDR;
input  [31:0] DW1;
input  [31:0] DW6;
input  [31:0] DW12;
input  [31:0] DW13;
output [3:0] SIDWOFFSET;
output [3:0] SIDWNUM;
input  [31:0] DW2;
input  [31:0] DW3;
input  [31:0] DW8;
input  [3:0] DWCNT;
output [13:0] SITDSM;
input  [31:0] DW4;
output [31:0] UP_DW5;
input  [10:0] ACTLEN;
input  [31:0] DW5;
input  [31:0] DW10;
input  [31:0] DW11;
output [31:0] UP_DW4;
output [104:0] TRAN_CMD;
output [31:0] UP_DW3;
input  SITD_PARSE_GO, GEN_PERR, PCIEND, SITD_ACT, CRCERR, BABBLE, PIDERR, 
    TMOUT, RXDATA0, RXDATA1, RXMDATA, RXNYET, RXPIDERR, EHCI_MAC_EOT, FEMPTY, 
    TDMAEND, SICMDSTART, HCI_PRESOF, LTINT_PCLK, USBINT_EN, ERRINT_EN, USBINT, 
    ERRINT, RECOVERYMODE, PCICLK, EHCIFLOW_PCLK, TRST_;
output PARSESITDEND, SITDPARSING, SITDIDLE, CACHEPHASE, UP_LDW3, UP_LDW4, 
    UP_LDW5, SIHCIREQ, SIHCIMWR, SIBUI_GO, CACHE_INVALID, SIRXERR, 
    SICMDSTART_REQ, SIEOT, SITDIOCINT_S, SITDERRINT_S, SITDIOCINT;
    wire SITDSMNXT_2, VIR_TOTALBYTES_9, TOTALBYTES621_2, CPROGMASK_COM_2, 
        NDW3_2, SIRXERR_CUR1009, SPAREO6, NDW3_25, HCI_PRESOF_T, TP757_1, 
        NDW3_19, RETRYCNT_0, OVERWBOFFSET_P1150_9, SMASK_2, IMMEDRETRY1046, 
        CMASK_1, VIR_TOTALBYTES_0, OVERWBOFFSET1181_6, OVERWBOFFSET1181_11, 
        SITDSMNXT_11, OVERWBOFFSET_P1150_0, RETRYCNT1099_1, CPROGMASK875_7, 
        NDW5_1, NDW3_30, NDW3_17, SITDIOCINT_T, CPROGMASK875_0, SPAREO0_, 
        OVERWBOFFSET_P1150_7, SPAREO8, OVERWBOFFSET1181_1, VIR_TOTALBYTES_7, 
        PG747, RETRYCNT1095_1, SMASK_5, CMASK_6, TCOUNT797_2, 
        OVERWBOFFSET_P1150_11, OVERWBOFFSET1181_8, NDW3_22, SPAREO1, 
        SITDSMNXT_5, CPROGMASK_COM_5, TOTALBYTES621_5, VIR_TOTALBYTES_6, 
        RETRYCNT1095_0, SPAREO9, OVERWBOFFSET1181_0, NDW3_16, CPROGMASK875_1, 
        PHASENXT_idle, OVERWBOFFSET_P1150_6, IMMEDRETRY, SPLITSTS, SITDSMNXT_4, 
        CPROGMASK_COM_4, NDW3_4, TOTALBYTES621_4, MISUF851, OVERWBOFFSET1181_9, 
        NDW3_23, SPAREO0, OVERWBOFFSET_P1150_10, SMASK_4, SPLITXSTATE_COM, 
        CMASK_7, SMASK_3, OVERWBOFFSET_12, CMASK_0, SITDERRINT_T, TP757_0, 
        NDW3_18, RETRYCNT_1, OVERWBOFFSET_P1150_8, TCOUNT793_2, SPLITXSTATE861, 
        SPAREO7, NDW3_24, SITDSMNXT_3, VIR_TOTALBYTES_8, TOTALBYTES621_3, 
        CPROGMASK_COM_3, NDW5_0, ACTIVE_COM, OVERWBOFFSET_P1150_1, 
        SITDSMNXT_10, CPROGMASK875_6, UP_CACHE1324, SITDIOCINT_T1478, 
        OVERWBOFFSET1181_7, OVERWBOFFSET1181_10, VIR_TOTALBYTES_1, ERR_STS831, 
        CPROGMASK_COM_1, TOTALBYTES621_1, CACHE_INVALID452, SIEOT1441, SPAREO5, 
        TCOUNT793_0, SICMDSTART_EOT, CMASK_2, LENGTMAX, SMASK_1, 
        TOTALBYTES621_8, BABBLE_STS841, SITDSMNXT_8, VIR_TOTALBYTES_3, 
        OVERWBOFFSET1181_5, OVERWBOFFSET1181_12, SICMDSTART_P, CPROGMASK875_4, 
        SITDSMNXT_12, OVERWBOFFSET_P1150_3, SPLITSTS1254, NDW5_2, 
        SITDERRINT_T1552, OVERWBOFFSET_P1150_4, CPROGMASK875_3, 
        PARSESITDEND_PRE, OVERWBOFFSET1181_2, VIR_TOTALBYTES_4, CMASK_5, 
        SMASK_6, OVERWBOFFSET_P1150_12, TCOUNT797_1, ACTIVE821, SPAREO2, 
        NDW3_21, BACKSTATE526, TOTALBYTES621_6, CPROGMASK_COM_6, NDW3_6, 
        SITDSMNXT_6, VIR_TOTALBYTES_5, SITDIOCINT1515, OVERWBOFFSET1181_3, 
        OVERWBOFFSET_P1150_5, CPROGMASK875_2, HCI_PRESOF_T489, NDW5_4, 
        TOTALBYTES621_7, CPROGMASK_COM_7, SITDSMNXT_7, SPAREO3, NDW3_20, 
        SPAREO1_, CMASK_4, UNDERFLOW, SMASK_7, CMASK_3, SMASK_0, n2176, 
        SPAREO4, TCOUNT793_1, CPROGMASK_COM_0, TOTALBYTES621_0, NDW5_3, 
        SICMDSTART_EOT1404, CPROGMASK875_5, OVERWBOFFSET_P1150_2, SITDSMNXT_13, 
        OVERWBOFFSET1181_4, TOTALBYTES621_9, SITDSMNXT_9, VIR_TOTALBYTES_2, 
        n1613, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, 
        n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, 
        n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, 
        n1775, n1779, n1781, n1782, n1783, n1784, n1815, n1816, n1817, n1818, 
        n1819, n1820, n1821, sub_342_carry_8, sub_342_carry_1, 
        sub_342_B_not_10, sub_342_B_not_8, sub_342_B_not_6, sub_342_B_not_1, 
        sub_342_carry_9, sub_342_carry_7, sub_342_carry_6, sub_342_B_not_7, 
        sub_342_B_not_9, sub_342_B_not_0, sub_342_carry_2, sub_342_B_not_5, 
        sub_342_B_not_2, sub_342_carry_10, sub_342_carry_5, sub_342_carry_4, 
        sub_342_B_not_4, sub_342_carry_3, sub_342_B_not_3, n1822, n1823, 
        r203_carry_8, r203_carry_1, r203_carry_12, r203_carry_7, r203_carry_6, 
        r203_carry_9, r203_carry_2, r203_carry_11, r203_carry_10, r203_carry_5, 
        r203_carry_4, r203_carry_3, n1824, n1825, n1826, n1827, n1828, n1829, 
        n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
        n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
        n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
        n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
        n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
        n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
        n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
        n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
        n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
        n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
        n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
        n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
        n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, 
        n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, 
        n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, 
        n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, 
        n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, 
        n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, 
        n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, 
        n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, 
        n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, 
        n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, 
        n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, 
        n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, 
        n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, 
        n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, 
        n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, 
        n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, 
        n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, 
        n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
        n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, 
        n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, 
        n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, 
        n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, 
        n2170, n2171, n2172, n2173, _cell_952_U2_Z_10, _cell_952_U2_Z_9, 
        _cell_952_U2_Z_8, _cell_952_U2_Z_7, _cell_952_U2_Z_6, _cell_952_U2_Z_5, 
        _cell_952_U2_Z_4, _cell_952_U2_Z_3, _cell_952_U2_Z_2, _cell_952_U2_Z_1, 
        _cell_952_U2_Z_0;
    assign UP_DW3[5] = 1'b0;
    assign SIDWNUM[3] = 1'b0;
    assign SIDWNUM[0] = 1'b0;
    assign SIDWOFFSET[3] = 1'b0;
    assign TRAN_CMD[51] = 1'b0;
    assign TRAN_CMD[50] = 1'b0;
    assign TRAN_CMD[11] = 1'b0;
    assign TRAN_CMD[10] = 1'b1;
    assign TRAN_CMD[7] = 1'b0;
    assign TRAN_CMD[6] = 1'b1;
    assign TRAN_CMD[5] = 1'b0;
    assign TRAN_CMD[4] = 1'b1;
    assign TRAN_CMD[2] = 1'b0;
    assign TRAN_CMD[0] = 1'b1;
    znd3b SPARE589 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE580 ( .CK(PCICLK), .D(IMMEDRETRY), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE587 ( .A(SPAREO4), .Y(SPAREO5) );
    znr3b SPARE586 ( .A(SPAREO2), .B(LENGTMAX), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE588 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE581 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zaoi211b SPARE583 ( .A(SPAREO4), .B(PARSESITDEND_PRE), .C(SPAREO6), .D(
        1'b0), .Y(SPAREO8) );
    zoai21b SPARE584 ( .A(SPAREO0), .B(SPAREO8), .C(n1751), .Y(SPAREO9) );
    zoai21b SPARE585 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE582 ( .A(SPAREO0), .B(n1773), .C(SPAREO1_), .D(SICMDSTART_P), 
        .Y(SPAREO2) );
    zxo2b U494 ( .A(n2075), .B(n1875), .Y(n2114) );
    zxo2b U495 ( .A(n2076), .B(n1874), .Y(n2113) );
    zxo2b U496 ( .A(n2074), .B(n1879), .Y(n2112) );
    zxo2b U497 ( .A(n2104), .B(n1876), .Y(n2111) );
    zxo2b U498 ( .A(n2071), .B(n1880), .Y(n2110) );
    zxo2b U499 ( .A(n2105), .B(n1877), .Y(n2109) );
    zxo2b U500 ( .A(CMASK_4), .B(n2128), .Y(n2108) );
    zxo2b U501 ( .A(n2072), .B(n1881), .Y(n2107) );
    zmux21lb U502 ( .A(n2064), .B(n2071), .S(n1752), .Y(n2134) );
    zmux21lb U503 ( .A(n2066), .B(n2073), .S(n1752), .Y(n2139) );
    zmux21lb U504 ( .A(n2068), .B(n2074), .S(n1752), .Y(n2136) );
    zmux21lb U505 ( .A(n2137), .B(n2105), .S(n1752), .Y(n2141) );
    zivb U506 ( .A(CMASK_4), .Y(n2073) );
    zivb U507 ( .A(CMASK_5), .Y(n2074) );
    zivb U508 ( .A(CMASK_6), .Y(n2071) );
    zivb U509 ( .A(SMASK_4), .Y(n2066) );
    zivb U510 ( .A(SMASK_5), .Y(n2068) );
    zivb U511 ( .A(SMASK_6), .Y(n2064) );
    zmux21lb U512 ( .A(SMASK_2), .B(CMASK_2), .S(n1752), .Y(n2129) );
    zmux21lb U513 ( .A(SMASK_1), .B(CMASK_1), .S(n1752), .Y(n2130) );
    znr3b U514 ( .A(n1816), .B(n1818), .C(n1815), .Y(n1817) );
    znd2b U515 ( .A(UP_DW3[19]), .B(UP_DW3[20]), .Y(n1816) );
    znr2b U516 ( .A(UP_DW3[16]), .B(UP_DW3[17]), .Y(n1818) );
    znd2b U517 ( .A(UP_DW3[18]), .B(UP_DW3[21]), .Y(n1815) );
    zan2b U518 ( .A(n1928), .B(n1929), .Y(n1927) );
    zao22b U519 ( .A(IMMEDRETRY), .B(n1841), .C(RXNYET), .D(n2162), .Y(n1995)
         );
    zivb U520 ( .A(n2106), .Y(n2162) );
    znd8b U521 ( .A(n2107), .B(n2108), .C(n2109), .D(n2110), .E(n2111), .F(
        n2112), .G(n2113), .H(n2114), .Y(n2106) );
    zoai2x4b U522 ( .A(n1926), .B(n2076), .C(n1925), .D(n2075), .E(n1913), .F(
        n2069), .G(n2062), .H(n2143), .Y(n1999) );
    zivb U523 ( .A(CMASK_1), .Y(n2075) );
    zmux21lb U524 ( .A(CMASK_2), .B(CMASK_3), .S(FRNUM[0]), .Y(n2143) );
    zivb U525 ( .A(CMASK_2), .Y(n2104) );
    zivb U526 ( .A(CMASK_3), .Y(n2105) );
    zoai2x4b U527 ( .A(n1926), .B(n1933), .C(n2070), .D(n1925), .E(n1917), .F(
        n2069), .G(n2062), .H(n2142), .Y(n1998) );
    zmux21lb U528 ( .A(SMASK_2), .B(SMASK_3), .S(FRNUM[0]), .Y(n2142) );
    zmux41b U529 ( .A(FRNUM[1]), .B(FRNUM[0]), .D0(n2140), .D1(n2135), .D2(
        n2138), .D3(n2133), .Y(n2082) );
    zan2b U530 ( .A(n2141), .B(n2127), .Y(n2140) );
    zan2b U531 ( .A(n2136), .B(n2125), .Y(n2135) );
    zan2b U532 ( .A(n2139), .B(n2126), .Y(n2138) );
    zan2b U533 ( .A(n2134), .B(n2124), .Y(n2133) );
    zan2b U534 ( .A(n1919), .B(n1920), .Y(n1918) );
    zmux21lb U535 ( .A(n2065), .B(n2072), .S(n1752), .Y(n1919) );
    zivb U536 ( .A(SMASK_7), .Y(n2065) );
    zivb U537 ( .A(CMASK_7), .Y(n2072) );
    zmux21lb U538 ( .A(n2131), .B(n2132), .S(FRNUM[0]), .Y(n2081) );
    zor2b U539 ( .A(CPROGMASK_COM_1), .B(n2130), .Y(n2131) );
    zor2b U540 ( .A(CPROGMASK_COM_2), .B(n2129), .Y(n2132) );
    zan2b U541 ( .A(n1922), .B(n1923), .Y(n1921) );
    zmux21lb U542 ( .A(n1933), .B(n2076), .S(n1752), .Y(n1922) );
    zivb U543 ( .A(CMASK_0), .Y(n2076) );
    znd2b U544 ( .A(UP_DW3[23]), .B(n1774), .Y(n1819) );
    znr2b U545 ( .A(UP_DW3[24]), .B(UP_DW3[25]), .Y(n1820) );
    zivb U546 ( .A(SMASK_0), .Y(n1933) );
    zivb U547 ( .A(SMASK_1), .Y(n2070) );
    zivb U548 ( .A(SMASK_3), .Y(n2137) );
    zoai2x4b U549 ( .A(n1958), .B(n2103), .C(n2158), .D(n2059), .E(n2000), .F(
        n2102), .G(n1959), .H(n1960), .Y(n2149) );
    zan2b U550 ( .A(n1959), .B(n1960), .Y(n1958) );
    zoai2x4b U551 ( .A(n1962), .B(n1963), .C(n1961), .D(n2083), .E(n2057), .F(
        n1977), .G(n2159), .H(n2160), .Y(n2147) );
    zan2b U552 ( .A(n1962), .B(n1963), .Y(n1961) );
    zivb U553 ( .A(n2048), .Y(n2160) );
    zan2b U554 ( .A(n1852), .B(n1980), .Y(n1979) );
    zxo2b U555 ( .A(n1821), .B(RETRYCNT_0), .Y(RETRYCNT1099_1) );
    zao21b U556 ( .A(n1821), .B(n2119), .C(n1772), .Y(n1994) );
    zoa211b U557 ( .A(SITDSM[9]), .B(SITDSM[7]), .C(SITD_ACT), .D(EHCI_MAC_EOT
        ), .Y(n2161) );
    zivb U558 ( .A(n1941), .Y(n1835) );
    zivb U559 ( .A(RXMDATA), .Y(n1991) );
    zcx4b U560 ( .A(n1930), .B(n1936), .C(n1937), .D(n1938), .Y(n1935) );
    zoa22b U561 ( .A(n1927), .B(n1931), .C(SPLITXSTATE_COM), .D(n1928), .Y(
        n1930) );
    zao22b U562 ( .A(n1756), .B(n1910), .C(FEMPTY), .D(n1760), .Y(n1938) );
    zivb U563 ( .A(ACTLEN[10]), .Y(sub_342_B_not_10) );
    znr2b U564 ( .A(UP_DW5[0]), .B(UP_DW5[1]), .Y(n1823) );
    zan3b U565 ( .A(n1822), .B(n1944), .C(n1945), .Y(n1943) );
    zor2b U566 ( .A(FRNUM[0]), .B(n2060), .Y(n2063) );
    zor2b U567 ( .A(FRNUM[1]), .B(FRNUM[0]), .Y(n2053) );
    zor2b U568 ( .A(FRNUM[2]), .B(n2060), .Y(n2062) );
    zivb U569 ( .A(FRNUM[1]), .Y(n2060) );
    zor2b U570 ( .A(FRNUM[1]), .B(n2061), .Y(n2067) );
    zivb U571 ( .A(n2067), .Y(n1916) );
    zor2b U572 ( .A(TRAN_CMD[8]), .B(n1940), .Y(n2086) );
    zan3b U573 ( .A(UP_DW3[1]), .B(n1941), .C(n1942), .Y(n1940) );
    zcx8d U574 ( .A(n1951), .B(n1928), .C(n1953), .D(n1954), .E(PCIEND), .Y(
        n1952) );
    zan2b U575 ( .A(UP_DW3[7]), .B(UP_DW3[1]), .Y(n2144) );
    znr8b U576 ( .A(n1990), .B(n1993), .C(n1994), .D(n1995), .E(RXDATA0), .F(
        RXDATA1), .G(RXPIDERR), .H(BABBLE), .Y(n1992) );
    zoa211b U577 ( .A(n1947), .B(n1950), .C(n1951), .D(n1931), .Y(n1949) );
    zan2b U578 ( .A(n1948), .B(SPLITXSTATE_COM), .Y(n1947) );
    zivb U579 ( .A(n1928), .Y(n1948) );
    zivb U580 ( .A(n1929), .Y(n1950) );
    zivb U581 ( .A(n1936), .Y(n1951) );
    zor2b U582 ( .A(n1997), .B(n2078), .Y(n1936) );
    zivb U583 ( .A(n1956), .Y(n2156) );
    zan2b U584 ( .A(SMASK_0), .B(n1754), .Y(n2154) );
    zor2b U585 ( .A(FRNUM[2]), .B(n2053), .Y(n1926) );
    zor2b U586 ( .A(SITDSM[12]), .B(SITDSM[9]), .Y(n2046) );
    zivb U587 ( .A(n2046), .Y(n2158) );
    zor2b U588 ( .A(SITDSM[10]), .B(n2046), .Y(n2047) );
    zivb U589 ( .A(n2047), .Y(n1959) );
    zoai2x4b U590 ( .A(n1921), .B(n1925), .C(n2062), .D(n2081), .E(n1918), .F(
        n1926), .G(n2069), .H(n2082), .Y(n1931) );
    zivb U591 ( .A(FRNUM[2]), .Y(n2069) );
    zmux21lb U592 ( .A(n1998), .B(n1999), .S(SPLITXSTATE_COM), .Y(n1997) );
    zor2b U593 ( .A(SITDSM[4]), .B(n2085), .Y(n1946) );
    zor2b U594 ( .A(SIDWOFFSET[2]), .B(n1868), .Y(n2152) );
    zor2b U595 ( .A(PARSESITDEND), .B(n1882), .Y(n2151) );
    zivb U596 ( .A(n2099), .Y(n2155) );
    zivb U597 ( .A(n2049), .Y(n2159) );
    zcx7b U598 ( .A(UP_DW3[1]), .B(TDMAEND), .C(n1975), .D(n1977), .E(n1978), 
        .Y(n1829) );
    znr8b U599 ( .A(n1976), .B(n1749), .C(n1750), .D(n1864), .E(n1863), .F(
        n1865), .G(n1867), .H(n1866), .Y(n1975) );
    znd2b U600 ( .A(n1820), .B(n1819), .Y(LENGTMAX) );
    zor2b U601 ( .A(TRAN_CMD[8]), .B(SPLITSTS), .Y(n1974) );
    zan2b U602 ( .A(n1966), .B(n1967), .Y(n1828) );
    zmux21hb U603 ( .A(n2050), .B(n2146), .S(n2150), .Y(n1826) );
    zor2b U604 ( .A(n2048), .B(n2049), .Y(n2050) );
    zivb U605 ( .A(n2050), .Y(n2148) );
    zivb U606 ( .A(n2055), .Y(n2150) );
    zor2b U607 ( .A(SIDWNUM[2]), .B(n2054), .Y(n2055) );
    zivb U608 ( .A(n1957), .Y(n1954) );
    zor2b U609 ( .A(UP_DW3[7]), .B(n1838), .Y(n1964) );
    zivb U610 ( .A(n1964), .Y(n1953) );
    zxo2b U611 ( .A(n1822), .B(UP_DW5[0]), .Y(TCOUNT797_1) );
    znd2b U612 ( .A(n1850), .B(n1851), .Y(RETRYCNT1095_1) );
    zmux21lb U613 ( .A(RETRYCNT_1), .B(RETRYCNT1099_1), .S(n1979), .Y(n1850)
         );
    zao32b U614 ( .A(n1852), .B(n2119), .C(n1853), .D(RETRYCNT_0), .E(n1854), 
        .Y(RETRYCNT1095_0) );
    zivb U615 ( .A(n2120), .Y(n1852) );
    zoai21b U616 ( .A(n1852), .B(n1861), .C(n2123), .Y(n1854) );
    zoai21b U617 ( .A(n1869), .B(n1870), .C(n1871), .Y(PG747) );
    zor2b U618 ( .A(n1981), .B(n1885), .Y(n1869) );
    zan2b U619 ( .A(SIDWOFFSET[2]), .B(n1984), .Y(n1857) );
    zivb U620 ( .A(n1969), .Y(SITDSMNXT_13) );
    zan2b U621 ( .A(SITDSM[12]), .B(n1838), .Y(UP_CACHE1324) );
    zao21b U622 ( .A(n2165), .B(n2161), .C(SIRXERR), .Y(n1899) );
    zivb U623 ( .A(n1899), .Y(n2121) );
    zivb U624 ( .A(n2085), .Y(SITDSMNXT_12) );
    zivb U625 ( .A(ACTLEN[9]), .Y(sub_342_B_not_9) );
    zivb U626 ( .A(VIR_TOTALBYTES_9), .Y(n1989) );
    zivb U627 ( .A(ACTLEN[8]), .Y(sub_342_B_not_8) );
    zivb U628 ( .A(VIR_TOTALBYTES_8), .Y(n1986) );
    zivb U629 ( .A(ACTLEN[7]), .Y(sub_342_B_not_7) );
    zivb U630 ( .A(VIR_TOTALBYTES_7), .Y(n2087) );
    zivb U631 ( .A(ACTLEN[6]), .Y(sub_342_B_not_6) );
    zivb U632 ( .A(VIR_TOTALBYTES_6), .Y(n2088) );
    zivb U633 ( .A(ACTLEN[5]), .Y(sub_342_B_not_5) );
    zivb U634 ( .A(VIR_TOTALBYTES_5), .Y(n2089) );
    zivb U635 ( .A(ACTLEN[4]), .Y(sub_342_B_not_4) );
    zivb U636 ( .A(VIR_TOTALBYTES_4), .Y(n2090) );
    zivb U637 ( .A(ACTLEN[3]), .Y(sub_342_B_not_3) );
    zivb U638 ( .A(VIR_TOTALBYTES_3), .Y(n2091) );
    zivb U639 ( .A(ACTLEN[2]), .Y(sub_342_B_not_2) );
    zivb U640 ( .A(VIR_TOTALBYTES_2), .Y(n2092) );
    zivb U641 ( .A(ACTLEN[1]), .Y(sub_342_B_not_1) );
    zivb U642 ( .A(VIR_TOTALBYTES_1), .Y(n2093) );
    zivb U643 ( .A(ACTLEN[0]), .Y(sub_342_B_not_0) );
    zivb U644 ( .A(VIR_TOTALBYTES_0), .Y(n2094) );
    zor2b U645 ( .A(n1939), .B(n1903), .Y(n1890) );
    zivb U646 ( .A(n2096), .Y(n2095) );
    zxo2b U647 ( .A(UP_DW5[2]), .B(n1823), .Y(TCOUNT797_2) );
    zao21b U648 ( .A(FRNUM[2]), .B(n1769), .C(UP_DW3[15]), .Y(n1881) );
    zao21b U649 ( .A(FRNUM[2]), .B(n1914), .C(UP_DW3[14]), .Y(n1880) );
    zivb U650 ( .A(n2063), .Y(n1914) );
    zao21b U651 ( .A(FRNUM[2]), .B(n1916), .C(UP_DW3[13]), .Y(n1879) );
    zao21b U652 ( .A(FRNUM[2]), .B(n1915), .C(UP_DW3[12]), .Y(n1878) );
    zivb U653 ( .A(n2053), .Y(n1915) );
    zivb U654 ( .A(CPROGMASK_COM_4), .Y(n2126) );
    zivb U655 ( .A(CPROGMASK_COM_5), .Y(n2125) );
    zivb U656 ( .A(CPROGMASK_COM_6), .Y(n2124) );
    zivb U657 ( .A(CPROGMASK_COM_7), .Y(n1920) );
    zivb U658 ( .A(n1878), .Y(n2128) );
    zao21b U659 ( .A(n2164), .B(FRNUM[0]), .C(UP_DW3[11]), .Y(n1877) );
    zao21b U660 ( .A(n2164), .B(n2061), .C(UP_DW3[10]), .Y(n1876) );
    zivb U661 ( .A(n2062), .Y(n2164) );
    zivb U662 ( .A(FRNUM[0]), .Y(n2061) );
    zor2b U663 ( .A(n2163), .B(UP_DW3[9]), .Y(n1875) );
    zivb U664 ( .A(n1925), .Y(n2163) );
    zor2b U665 ( .A(n1982), .B(n1903), .Y(n1872) );
    zao21b U666 ( .A(UP_DW3[1]), .B(n1853), .C(n1765), .Y(n1873) );
    zor2b U667 ( .A(n2157), .B(UP_DW3[8]), .Y(n1874) );
    zivb U668 ( .A(n1926), .Y(n2157) );
    zivb U669 ( .A(CPROGMASK_COM_0), .Y(n1923) );
    zivb U670 ( .A(CPROGMASK_COM_3), .Y(n2127) );
    zao22b U671 ( .A(n1906), .B(n1853), .C(OVERWBOFFSET_12), .D(n1903), .Y(
        OVERWBOFFSET1181_12) );
    zivb U672 ( .A(n1870), .Y(n1906) );
    znd2b U673 ( .A(OVERWBOFFSET_P1150_12), .B(n2086), .Y(n1870) );
    zivd U674 ( .A(n2123), .Y(n1903) );
    zor2b U675 ( .A(n1980), .B(n1861), .Y(n2123) );
    zivc U676 ( .A(n2122), .Y(n1904) );
    zor2b U677 ( .A(n1981), .B(n1885), .Y(n2122) );
    zivb U678 ( .A(n2086), .Y(n1981) );
    zan2b U679 ( .A(n1841), .B(n1868), .Y(HCI_PRESOF_T489) );
    zivb U680 ( .A(n1858), .Y(SITDSMNXT_3) );
    zmux31hb U681 ( .A(n1851), .B(SITDSM[3]), .D0(SPLITXSTATE_COM), .D1(UP_DW3
        [1]), .D2(n2144), .Y(n1884) );
    zivb U682 ( .A(n1965), .Y(n1908) );
    zor2b U683 ( .A(SITDSM[4]), .B(SITDSM[2]), .Y(n1965) );
    zivb U684 ( .A(n2051), .Y(n1909) );
    zmux21lb U685 ( .A(n2078), .B(n2153), .S(n1851), .Y(ACTIVE821) );
    zor2b U686 ( .A(n1751), .B(n1839), .Y(n2153) );
    zmux21lb U687 ( .A(n2077), .B(n2145), .S(n1851), .Y(SPLITSTS1254) );
    zivb U688 ( .A(SPLITXSTATE_COM), .Y(n2077) );
    zmux21lb U689 ( .A(SPLITSTS), .B(UP_DW3[1]), .S(SIBUI_GO), .Y(n2145) );
    zivb U690 ( .A(n2100), .Y(SITDSMNXT_5) );
    zoai21b U691 ( .A(n2101), .B(n1949), .C(n1832), .Y(n2100) );
    zoai21b U692 ( .A(n1885), .B(n1886), .C(n1887), .Y(BABBLE_STS841) );
    zivb U693 ( .A(BABBLE), .Y(n1886) );
    zmux21lb U694 ( .A(NDW3_4), .B(UP_DW3[4]), .S(n1851), .Y(n1887) );
    zoai21b U695 ( .A(n1885), .B(n1896), .C(n1897), .Y(ERR_STS831) );
    zor2b U696 ( .A(n1946), .B(n1861), .Y(n1885) );
    zmux21lb U697 ( .A(NDW3_6), .B(UP_DW3[6]), .S(n1851), .Y(n1897) );
    zivb U698 ( .A(n1885), .Y(n1853) );
    zan3b U699 ( .A(n1882), .B(n1868), .C(n1883), .Y(IMMEDRETRY1046) );
    zivb U700 ( .A(SITD_PARSE_GO), .Y(n1882) );
    zmux21lb U701 ( .A(n2098), .B(n2120), .S(n1980), .Y(n1883) );
    zivb U702 ( .A(n1946), .Y(n1980) );
    zoa211b U703 ( .A(SITDIOCINT), .B(n1901), .C(n1902), .D(USBINT_EN), .Y(
        SITDIOCINT1515) );
    znd2b U704 ( .A(USBINT), .B(LTINT_PCLK), .Y(n1902) );
    zan2b U705 ( .A(n1911), .B(n1832), .Y(SITDSMNXT_11) );
    zao22b U706 ( .A(n1760), .B(n2084), .C(n1942), .D(n1759), .Y(n1911) );
    zivb U707 ( .A(FEMPTY), .Y(n2084) );
    zao33b U708 ( .A(n1758), .B(n1832), .C(n1833), .D(n1757), .E(SICMDSTART), 
        .F(n1764), .Y(SITDSMNXT_9) );
    zmux21hb U709 ( .A(NDW3_2), .B(n1993), .S(n1851), .Y(MISUF851) );
    zor2b U710 ( .A(UP_DW3[2]), .B(n1773), .Y(n1993) );
    zivb U711 ( .A(ACTIVE_COM), .Y(n2078) );
    zor2b U712 ( .A(SITDSM[6]), .B(SITDSM[8]), .Y(n1840) );
    zor2b U713 ( .A(HCI_PRESOF), .B(HCI_PRESOF_T), .Y(n1841) );
    zan2b U714 ( .A(n1910), .B(SITDSM[7]), .Y(n1842) );
    zivb U715 ( .A(n1840), .Y(n1962) );
    zao33b U716 ( .A(n1756), .B(n1832), .C(n1833), .D(SICMDSTART), .E(n1755), 
        .F(n1764), .Y(SITDSMNXT_7) );
    zivb U717 ( .A(SITDSMNXT_7), .Y(n1978) );
    zmux21lb U718 ( .A(n2151), .B(n2152), .S(n1837), .Y(n1844) );
    zoai21b U719 ( .A(LTINT_PCLK), .B(n1855), .C(n1856), .Y(SITDIOCINT_T1478)
         );
    zivb U720 ( .A(n1901), .Y(n1856) );
    zor2b U721 ( .A(SIRXERR), .B(BABBLE), .Y(n1888) );
    zan2b U722 ( .A(SITDERRINT_T), .B(n1970), .Y(n1889) );
    zivb U723 ( .A(LTINT_PCLK), .Y(n1970) );
    zivb U724 ( .A(n1888), .Y(n1942) );
    zao32b U725 ( .A(n1755), .B(n1898), .C(n1764), .D(n1766), .E(n1847), .Y(
        SITDSMNXT_6) );
    zan3b U726 ( .A(n1758), .B(n1832), .C(n1910), .Y(SITDSMNXT_10) );
    zivb U727 ( .A(n1833), .Y(n1910) );
    zor2b U728 ( .A(SICMDSTART), .B(n1845), .Y(n1833) );
    zao32b U729 ( .A(n1757), .B(n1898), .C(n1764), .D(n1766), .E(TRAN_CMD[104]
        ), .Y(SITDSMNXT_8) );
    zivb U730 ( .A(SICMDSTART), .Y(n1898) );
    zivb U731 ( .A(EHCI_MAC_EOT), .Y(n1845) );
    zan2b U732 ( .A(SITDERRINT_T), .B(LTINT_PCLK), .Y(SITDERRINT_S) );
    zan2b U733 ( .A(LTINT_PCLK), .B(SITDIOCINT_T), .Y(SITDIOCINT_S) );
    zan2b U734 ( .A(SICMDSTART_P), .B(n1843), .Y(SICMDSTART_REQ) );
    zivb U735 ( .A(n1900), .Y(SIBUI_GO) );
    zor2b U736 ( .A(SITDSM[5]), .B(n2100), .Y(n1900) );
    zan2b U737 ( .A(n1849), .B(n1847), .Y(TRAN_CMD[12]) );
    zxo2b U738 ( .A(n1996), .B(UP_DW5[4]), .Y(n1849) );
    zivb U739 ( .A(n1849), .Y(n1892) );
    zan2b U740 ( .A(n1847), .B(n1848), .Y(TRAN_CMD[13]) );
    zan2b U741 ( .A(n1746), .B(n1862), .Y(TRAN_CMD[40]) );
    zan2b U742 ( .A(n1750), .B(n1862), .Y(TRAN_CMD[41]) );
    zan2b U743 ( .A(n1867), .B(n1862), .Y(TRAN_CMD[42]) );
    zor2b U744 ( .A(n1761), .B(UP_DW3[18]), .Y(n1867) );
    zan2b U745 ( .A(n1866), .B(n1862), .Y(TRAN_CMD[43]) );
    zor2b U746 ( .A(n1761), .B(UP_DW3[19]), .Y(n1866) );
    zan2b U747 ( .A(n1865), .B(n1862), .Y(TRAN_CMD[44]) );
    zor2b U748 ( .A(n1761), .B(UP_DW3[20]), .Y(n1865) );
    zan2b U749 ( .A(n1864), .B(n1862), .Y(TRAN_CMD[45]) );
    zor2b U750 ( .A(n1761), .B(UP_DW3[21]), .Y(n1864) );
    zan2b U751 ( .A(n1747), .B(n1862), .Y(TRAN_CMD[46]) );
    zan2b U752 ( .A(n1863), .B(n1862), .Y(TRAN_CMD[47]) );
    zor2b U753 ( .A(n1761), .B(UP_DW3[23]), .Y(n1863) );
    zan2b U754 ( .A(n1749), .B(n1862), .Y(TRAN_CMD[48]) );
    zan2b U755 ( .A(n1748), .B(n1862), .Y(TRAN_CMD[49]) );
    zivb U756 ( .A(TRAN_CMD[104]), .Y(n1847) );
    zivd U757 ( .A(n2118), .Y(n2167) );
    zivd U758 ( .A(n2117), .Y(n1895) );
    zivb U759 ( .A(DWCNT[0]), .Y(n2116) );
    zivd U760 ( .A(n2118), .Y(n1893) );
    zivd U761 ( .A(n2117), .Y(n2170) );
    zan2b U762 ( .A(DW6[0]), .B(SIDWOFFSET[2]), .Y(SIHCIADR[0]) );
    zan2b U763 ( .A(DW6[1]), .B(SIDWOFFSET[2]), .Y(SIHCIADR[1]) );
    zan2b U764 ( .A(DW6[4]), .B(n1860), .Y(SIHCIADR[4]) );
    zao22b U765 ( .A(CACHE_ADDR[0]), .B(n1859), .C(DW6[5]), .D(n1860), .Y(
        SIHCIADR[5]) );
    zao22b U766 ( .A(CACHE_ADDR[1]), .B(n2171), .C(DW6[6]), .D(n2172), .Y(
        SIHCIADR[6]) );
    zao22b U767 ( .A(CACHE_ADDR[2]), .B(n1859), .C(DW6[7]), .D(n2173), .Y(
        SIHCIADR[7]) );
    zao22b U768 ( .A(CACHE_ADDR[3]), .B(n2171), .C(DW6[8]), .D(n1860), .Y(
        SIHCIADR[8]) );
    zao22b U769 ( .A(n1859), .B(CACHE_ADDR[4]), .C(DW6[9]), .D(n2172), .Y(
        SIHCIADR[9]) );
    zao22b U770 ( .A(CACHE_ADDR[5]), .B(n1859), .C(DW6[10]), .D(n2173), .Y(
        SIHCIADR[10]) );
    zao22b U771 ( .A(CACHE_ADDR[6]), .B(n2171), .C(DW6[11]), .D(n1860), .Y(
        SIHCIADR[11]) );
    zao22b U772 ( .A(CACHE_ADDR[7]), .B(n1859), .C(DW6[12]), .D(n2173), .Y(
        SIHCIADR[12]) );
    zao22b U773 ( .A(CACHE_ADDR[8]), .B(n2171), .C(DW6[13]), .D(n2172), .Y(
        SIHCIADR[13]) );
    zao22b U774 ( .A(CACHE_ADDR[9]), .B(n1859), .C(DW6[14]), .D(n1860), .Y(
        SIHCIADR[14]) );
    zao22b U775 ( .A(CACHE_ADDR[10]), .B(n2171), .C(DW6[15]), .D(n2172), .Y(
        SIHCIADR[15]) );
    zao22b U776 ( .A(CACHE_ADDR[11]), .B(n1859), .C(DW6[16]), .D(n2173), .Y(
        SIHCIADR[16]) );
    zao22b U777 ( .A(CACHE_ADDR[12]), .B(n2171), .C(DW6[17]), .D(n1860), .Y(
        SIHCIADR[17]) );
    zao22b U778 ( .A(CACHE_ADDR[13]), .B(n1859), .C(DW6[18]), .D(n2173), .Y(
        SIHCIADR[18]) );
    zao22b U779 ( .A(CACHE_ADDR[14]), .B(n2171), .C(DW6[19]), .D(n2172), .Y(
        SIHCIADR[19]) );
    zao22b U780 ( .A(CACHE_ADDR[15]), .B(n1859), .C(DW6[20]), .D(n1860), .Y(
        SIHCIADR[20]) );
    zao22b U781 ( .A(CACHE_ADDR[16]), .B(n2171), .C(DW6[21]), .D(n2172), .Y(
        SIHCIADR[21]) );
    zao22b U782 ( .A(CACHE_ADDR[17]), .B(n1859), .C(DW6[22]), .D(n2173), .Y(
        SIHCIADR[22]) );
    zao22b U783 ( .A(CACHE_ADDR[18]), .B(n2171), .C(DW6[23]), .D(n1860), .Y(
        SIHCIADR[23]) );
    zao22b U784 ( .A(CACHE_ADDR[19]), .B(n1859), .C(DW6[24]), .D(n2172), .Y(
        SIHCIADR[24]) );
    zao22b U785 ( .A(CACHE_ADDR[20]), .B(n2171), .C(DW6[25]), .D(n2173), .Y(
        SIHCIADR[25]) );
    zao22b U786 ( .A(CACHE_ADDR[21]), .B(n1859), .C(DW6[26]), .D(n1860), .Y(
        SIHCIADR[26]) );
    zao22b U787 ( .A(CACHE_ADDR[22]), .B(n2171), .C(DW6[27]), .D(n2172), .Y(
        SIHCIADR[27]) );
    zao22b U788 ( .A(CACHE_ADDR[23]), .B(n1859), .C(DW6[28]), .D(n2173), .Y(
        SIHCIADR[28]) );
    zao22b U789 ( .A(CACHE_ADDR[24]), .B(n2171), .C(DW6[29]), .D(n1860), .Y(
        SIHCIADR[29]) );
    zao22b U790 ( .A(CACHE_ADDR[25]), .B(n1859), .C(DW6[30]), .D(n2172), .Y(
        SIHCIADR[30]) );
    zor2b U791 ( .A(SIDWOFFSET[2]), .B(n1753), .Y(n2172) );
    zao22b U792 ( .A(CACHE_ADDR[26]), .B(n2171), .C(DW6[31]), .D(n2173), .Y(
        SIHCIADR[31]) );
    zivc U793 ( .A(n2115), .Y(n2171) );
    zor2b U794 ( .A(SIDWOFFSET[2]), .B(n1784), .Y(n2115) );
    zor2b U795 ( .A(SIDWOFFSET[2]), .B(n1753), .Y(n2173) );
    zivd U796 ( .A(n2115), .Y(n1859) );
    zivb U797 ( .A(n2079), .Y(n1966) );
    zivb U798 ( .A(n1967), .Y(n1971) );
    zor2b U799 ( .A(n1846), .B(SIDWNUM[2]), .Y(SIDWNUM[1]) );
    zivb U800 ( .A(RXPIDERR), .Y(n1896) );
    zivb U801 ( .A(RXNYET), .Y(n1973) );
    zor2b U802 ( .A(SITDSM[13]), .B(SIDWNUM[2]), .Y(SIHCIREQ) );
    zivb U803 ( .A(UP_DW5[12]), .Y(n2031) );
    zivb U804 ( .A(UP_DW5[13]), .Y(n2029) );
    zivb U805 ( .A(UP_DW5[14]), .Y(n2027) );
    zivb U806 ( .A(UP_DW5[15]), .Y(n2025) );
    zivb U807 ( .A(UP_DW5[16]), .Y(n2023) );
    zivb U808 ( .A(UP_DW5[17]), .Y(n2021) );
    zivb U809 ( .A(UP_DW5[18]), .Y(n2019) );
    zivb U810 ( .A(UP_DW5[19]), .Y(n2017) );
    zivb U811 ( .A(UP_DW5[20]), .Y(n2015) );
    zivb U812 ( .A(UP_DW5[21]), .Y(n2013) );
    zivb U813 ( .A(UP_DW5[22]), .Y(n2011) );
    zivb U814 ( .A(UP_DW5[23]), .Y(n2009) );
    zivb U815 ( .A(UP_DW5[24]), .Y(n2007) );
    zivb U816 ( .A(UP_DW5[25]), .Y(n2005) );
    zivb U817 ( .A(UP_DW5[26]), .Y(n2003) );
    zivb U818 ( .A(UP_DW5[27]), .Y(n2001) );
    zivb U819 ( .A(UP_DW5[28]), .Y(n2044) );
    zivb U820 ( .A(UP_DW5[29]), .Y(n2042) );
    zivb U821 ( .A(UP_DW5[30]), .Y(n2040) );
    zivb U822 ( .A(UP_DW5[31]), .Y(n2038) );
    zivb U823 ( .A(UP_DW4[12]), .Y(n2032) );
    zivb U824 ( .A(UP_DW4[13]), .Y(n2030) );
    zivb U825 ( .A(UP_DW4[14]), .Y(n2028) );
    zivb U826 ( .A(UP_DW4[15]), .Y(n2026) );
    zivb U827 ( .A(UP_DW4[16]), .Y(n2024) );
    zivb U828 ( .A(UP_DW4[17]), .Y(n2022) );
    zivb U829 ( .A(UP_DW4[18]), .Y(n2020) );
    zivb U830 ( .A(UP_DW4[19]), .Y(n2018) );
    zivb U831 ( .A(UP_DW4[20]), .Y(n2016) );
    zivb U832 ( .A(UP_DW4[21]), .Y(n2014) );
    zivb U833 ( .A(UP_DW4[22]), .Y(n2012) );
    zivb U834 ( .A(UP_DW4[23]), .Y(n2010) );
    zivb U835 ( .A(UP_DW4[24]), .Y(n2008) );
    zivb U836 ( .A(UP_DW4[25]), .Y(n2006) );
    zivb U837 ( .A(UP_DW4[26]), .Y(n2004) );
    zivb U838 ( .A(UP_DW4[27]), .Y(n2002) );
    zivb U839 ( .A(UP_DW4[28]), .Y(n2045) );
    zivb U840 ( .A(UP_DW4[29]), .Y(n2043) );
    zivb U841 ( .A(UP_DW4[30]), .Y(n2041) );
    zivb U842 ( .A(UP_DW4[31]), .Y(n2039) );
    zan2b U843 ( .A(n1836), .B(n1837), .Y(SITDPARSING) );
    zivb U844 ( .A(PHASENXT_idle), .Y(n1837) );
    zivb U845 ( .A(SITDSM[13]), .Y(n2103) );
    zbfb U846 ( .A(UP_LDW3), .Y(UP_LDW5) );
    zivb U847 ( .A(SITDSM[12]), .Y(n2000) );
    zivb U848 ( .A(SITDSM[0]), .Y(n1868) );
    zdffqrb TOTALBYTES_reg_9 ( .CK(PCICLK), .D(TOTALBYTES621_9), .R(TRST_), 
        .Q(UP_DW3[25]) );
    zivb U849 ( .A(UP_DW3[25]), .Y(n2033) );
    zdffqrb TOTALBYTES_reg_8 ( .CK(PCICLK), .D(TOTALBYTES621_8), .R(TRST_), 
        .Q(UP_DW3[24]) );
    zivb U850 ( .A(UP_DW3[24]), .Y(n2034) );
    zdffqrb TOTALBYTES_reg_7 ( .CK(PCICLK), .D(TOTALBYTES621_7), .R(TRST_), 
        .Q(UP_DW3[23]) );
    zdffqrb TOTALBYTES_reg_6 ( .CK(PCICLK), .D(TOTALBYTES621_6), .R(TRST_), 
        .Q(UP_DW3[22]) );
    zivb U851 ( .A(UP_DW3[22]), .Y(n2035) );
    zdffqrb TOTALBYTES_reg_5 ( .CK(PCICLK), .D(TOTALBYTES621_5), .R(TRST_), 
        .Q(UP_DW3[21]) );
    zdffqrb TOTALBYTES_reg_4 ( .CK(PCICLK), .D(TOTALBYTES621_4), .R(TRST_), 
        .Q(UP_DW3[20]) );
    zdffqrb TOTALBYTES_reg_3 ( .CK(PCICLK), .D(TOTALBYTES621_3), .R(TRST_), 
        .Q(UP_DW3[19]) );
    zdffqrb TOTALBYTES_reg_2 ( .CK(PCICLK), .D(TOTALBYTES621_2), .R(TRST_), 
        .Q(UP_DW3[18]) );
    zdffqrb TOTALBYTES_reg_1 ( .CK(PCICLK), .D(TOTALBYTES621_1), .R(TRST_), 
        .Q(UP_DW3[17]) );
    zivb U852 ( .A(UP_DW3[17]), .Y(n2036) );
    zdffqrb TOTALBYTES_reg_0 ( .CK(PCICLK), .D(TOTALBYTES621_0), .R(TRST_), 
        .Q(UP_DW3[16]) );
    zivb U853 ( .A(UP_DW3[16]), .Y(n2037) );
    zdffqb TP_reg_1 ( .CK(PCICLK), .D(TP757_1), .Q(UP_DW5[4]) );
    zivb U854 ( .A(UP_DW5[4]), .Y(n1848) );
    zdffqb TP_reg_0 ( .CK(PCICLK), .D(TP757_0), .Q(UP_DW5[3]) );
    zivb U855 ( .A(UP_DW5[3]), .Y(n1996) );
    zdffqb TCOUNT_reg_2 ( .CK(PCICLK), .D(TCOUNT793_2), .Q(UP_DW5[2]) );
    zivb U856 ( .A(UP_DW5[2]), .Y(n1944) );
    zdffqb CPROGMASK_reg_7 ( .CK(PCICLK), .D(CPROGMASK875_7), .Q(UP_DW3[15])
         );
    zdffqb CPROGMASK_reg_6 ( .CK(PCICLK), .D(CPROGMASK875_6), .Q(UP_DW3[14])
         );
    zdffqb CPROGMASK_reg_5 ( .CK(PCICLK), .D(CPROGMASK875_5), .Q(UP_DW3[13])
         );
    zdffqb CPROGMASK_reg_4 ( .CK(PCICLK), .D(CPROGMASK875_4), .Q(UP_DW3[12])
         );
    zdffqb CPROGMASK_reg_3 ( .CK(PCICLK), .D(CPROGMASK875_3), .Q(UP_DW3[11])
         );
    zdffqb CPROGMASK_reg_2 ( .CK(PCICLK), .D(CPROGMASK875_2), .Q(UP_DW3[10])
         );
    zdffqb CPROGMASK_reg_1 ( .CK(PCICLK), .D(CPROGMASK875_1), .Q(UP_DW3[9]) );
    zdffqb CPROGMASK_reg_0 ( .CK(PCICLK), .D(CPROGMASK875_0), .Q(UP_DW3[8]) );
    zdffqb OVERWBOFFSET_reg_12 ( .CK(PCICLK), .D(OVERWBOFFSET1181_12), .Q(
        OVERWBOFFSET_12) );
    zdffqb OVERWBOFFSET_reg_11 ( .CK(PCICLK), .D(OVERWBOFFSET1181_11), .Q(
        UP_DW4[11]) );
    zdffqb OVERWBOFFSET_reg_10 ( .CK(PCICLK), .D(OVERWBOFFSET1181_10), .Q(
        UP_DW4[10]) );
    zdffqb OVERWBOFFSET_reg_9 ( .CK(PCICLK), .D(OVERWBOFFSET1181_9), .Q(UP_DW4
        [9]) );
    zdffqb OVERWBOFFSET_reg_8 ( .CK(PCICLK), .D(OVERWBOFFSET1181_8), .Q(UP_DW4
        [8]) );
    zdffqb OVERWBOFFSET_reg_7 ( .CK(PCICLK), .D(OVERWBOFFSET1181_7), .Q(UP_DW4
        [7]) );
    zdffqb OVERWBOFFSET_reg_6 ( .CK(PCICLK), .D(OVERWBOFFSET1181_6), .Q(UP_DW4
        [6]) );
    zdffqb OVERWBOFFSET_reg_5 ( .CK(PCICLK), .D(OVERWBOFFSET1181_5), .Q(UP_DW4
        [5]) );
    zdffqb OVERWBOFFSET_reg_4 ( .CK(PCICLK), .D(OVERWBOFFSET1181_4), .Q(UP_DW4
        [4]) );
    zdffqb OVERWBOFFSET_reg_3 ( .CK(PCICLK), .D(OVERWBOFFSET1181_3), .Q(UP_DW4
        [3]) );
    zdffqb OVERWBOFFSET_reg_2 ( .CK(PCICLK), .D(OVERWBOFFSET1181_2), .Q(UP_DW4
        [2]) );
    zdffqb OVERWBOFFSET_reg_1 ( .CK(PCICLK), .D(OVERWBOFFSET1181_1), .Q(UP_DW4
        [1]) );
    zdffqb OVERWBOFFSET_reg_0 ( .CK(PCICLK), .D(OVERWBOFFSET1181_0), .Q(UP_DW4
        [0]) );
    zdffqrb HCI_PRESOF_T_reg ( .CK(PCICLK), .D(HCI_PRESOF_T489), .R(TRST_), 
        .Q(HCI_PRESOF_T) );
    zdffqrb SITDSM_reg_3 ( .CK(PCICLK), .D(SITDSMNXT_3), .R(TRST_), .Q(SITDSM
        [3]) );
    zivb U857 ( .A(UP_DW3[1]), .Y(n1983) );
    zdffrb SITDSM_reg_4 ( .CK(PCICLK), .D(SITDSMNXT_4), .R(TRST_), .Q(SITDSM
        [4]), .QN(n2052) );
    zdffqrb SICMDSTART_EOT_reg ( .CK(PCICLK), .D(SICMDSTART_EOT1404), .R(TRST_
        ), .Q(SICMDSTART_EOT) );
    zivb U858 ( .A(SICMDSTART_EOT), .Y(n1843) );
    zdffqb ACTIVE_reg ( .CK(PCICLK), .D(ACTIVE821), .Q(UP_DW3[7]) );
    zivb U859 ( .A(UP_DW3[7]), .Y(n1839) );
    zdffqrb SPLITSTS_reg ( .CK(PCICLK), .D(SPLITSTS1254), .R(TRST_), .Q(
        SPLITSTS) );
    zdffqrb SITDSM_reg_5 ( .CK(PCICLK), .D(SITDSMNXT_5), .R(TRST_), .Q(SITDSM
        [5]) );
    zivb U860 ( .A(SITDSM[5]), .Y(n1963) );
    zdffqb BABBLE_STS_reg ( .CK(PCICLK), .D(BABBLE_STS841), .Q(UP_DW3[4]) );
    zdffqb ERR_STS_reg ( .CK(PCICLK), .D(ERR_STS831), .Q(UP_DW3[6]) );
    zdffqrb SITDSM_reg_2 ( .CK(PCICLK), .D(SITDSMNXT_2), .R(TRST_), .Q(SITDSM
        [2]) );
    zivb U861 ( .A(SITDSM[2]), .Y(n2080) );
    zdffqrb IMMEDRETRY_reg ( .CK(PCICLK), .D(IMMEDRETRY1046), .R(TRST_), .Q(
        IMMEDRETRY) );
    zivb U862 ( .A(IMMEDRETRY), .Y(n2098) );
    zdffqrb SITDIOCINT_reg ( .CK(EHCIFLOW_PCLK), .D(SITDIOCINT1515), .R(TRST_), 
        .Q(SITDIOCINT) );
    zdffqrb SITDSM_reg_11 ( .CK(PCICLK), .D(SITDSMNXT_11), .R(TRST_), .Q(
        SITDSM[11]) );
    zivb U863 ( .A(SITDSM[11]), .Y(n1960) );
    zdffqrb SITDSM_reg_9 ( .CK(PCICLK), .D(SITDSMNXT_9), .R(TRST_), .Q(SITDSM
        [9]) );
    zivb U864 ( .A(SITDSM[9]), .Y(n2102) );
    zdffqrb CACHE_INVALID_reg ( .CK(PCICLK), .D(CACHE_INVALID452), .R(TRST_), 
        .Q(CACHE_INVALID) );
    zdffqb MISUF_reg ( .CK(PCICLK), .D(MISUF851), .Q(UP_DW3[2]) );
    zivb U865 ( .A(UP_DW3[2]), .Y(n1972) );
    zdffqrb SIEOT_reg ( .CK(PCICLK), .D(SIEOT1441), .R(TRST_), .Q(SIEOT) );
    zdffqrb SITDSM_reg_7 ( .CK(PCICLK), .D(SITDSMNXT_7), .R(TRST_), .Q(SITDSM
        [7]) );
    zivb U866 ( .A(SITDSM[7]), .Y(n2083) );
    zdffqrb PARSESITDEND_reg ( .CK(PCICLK), .D(PARSESITDEND_PRE), .R(TRST_), 
        .Q(PARSESITDEND) );
    zdffqrb SITDIOCINT_T_reg ( .CK(EHCIFLOW_PCLK), .D(SITDIOCINT_T1478), .R(
        TRST_), .Q(SITDIOCINT_T) );
    zivb U867 ( .A(SITDIOCINT_T), .Y(n1855) );
    zdffqrb SITDERRINT_T_reg ( .CK(EHCIFLOW_PCLK), .D(SITDERRINT_T1552), .R(
        TRST_), .Q(SITDERRINT_T) );
    zdffqrb SITDSM_reg_6 ( .CK(PCICLK), .D(SITDSMNXT_6), .R(TRST_), .Q(SITDSM
        [6]) );
    zivb U868 ( .A(SITDSM[6]), .Y(n1977) );
    zdffqrb SITDSM_reg_10 ( .CK(PCICLK), .D(SITDSMNXT_10), .R(TRST_), .Q(
        SITDSM[10]) );
    zivb U869 ( .A(SITDSM[10]), .Y(n2059) );
    zdffqrb SITDSM_reg_8 ( .CK(PCICLK), .D(SITDSMNXT_8), .R(TRST_), .Q(SITDSM
        [8]) );
    zivb U870 ( .A(SITDSM[8]), .Y(n2057) );
    zivb U871 ( .A(SIDWNUM[2]), .Y(n1984) );
    zdffb TCOUNT_reg_1 ( .CK(PCICLK), .D(TCOUNT793_1), .Q(UP_DW5[1]), .QN(
        n1822) );
    znr2b U872 ( .A(n1761), .B(n2037), .Y(n1746) );
    znr2b U873 ( .A(n1761), .B(n2035), .Y(n1747) );
    znr2b U874 ( .A(n1761), .B(n2033), .Y(n1748) );
    znr2b U875 ( .A(n1761), .B(n2034), .Y(n1749) );
    zdffb RETRYCNT_reg_1 ( .CK(PCICLK), .D(RETRYCNT1095_1), .Q(RETRYCNT_1), 
        .QN(n1821) );
    znr2b U876 ( .A(n1761), .B(n2036), .Y(n1750) );
    znr2b U877 ( .A(n1992), .B(n1946), .Y(n1751) );
    znr2d U878 ( .A(TRAN_CMD[8]), .B(n2077), .Y(n1752) );
    znr2d U879 ( .A(SIDWOFFSET[2]), .B(n1838), .Y(n1753) );
    znr4b U880 ( .A(SITDSM[2]), .B(SITDSM[3]), .C(n2052), .D(n2051), .Y(n1754)
         );
    znr4b U881 ( .A(SITDSM[8]), .B(SITDSM[5]), .C(n1977), .D(n2056), .Y(n1755)
         );
    znr5b U882 ( .A(SITDSM[5]), .B(n1840), .C(n2049), .D(n2055), .E(n2083), 
        .Y(n1756) );
    znr4b U883 ( .A(SITDSM[6]), .B(SITDSM[5]), .C(n2057), .D(n2056), .Y(n1757)
         );
    znr3b U884 ( .A(SITDSM[12]), .B(n2102), .C(n2097), .Y(n1758) );
    znr4b U885 ( .A(SITDSM[11]), .B(n2046), .C(n2059), .D(n2058), .Y(n1759) );
    znr3b U886 ( .A(n2047), .B(n1960), .C(n2058), .Y(n1760) );
    zan2d U887 ( .A(LENGTMAX), .B(TRAN_CMD[8]), .Y(n1761) );
    znr2d U888 ( .A(UNDERFLOW), .B(n1869), .Y(n1762) );
    znr4b U889 ( .A(n2050), .B(n2054), .C(n1984), .D(GEN_PERR), .Y(n1763) );
    znr2b U890 ( .A(GEN_PERR), .B(n1841), .Y(n1764) );
    znr2b U891 ( .A(n2176), .B(n1885), .Y(n1765) );
    znr3b U892 ( .A(n2099), .B(n1845), .C(GEN_PERR), .Y(n1766) );
    znr2b U893 ( .A(n2166), .B(n2096), .Y(n1767) );
    znr2b U894 ( .A(n2095), .B(n2166), .Y(n1768) );
    znr2b U895 ( .A(n2060), .B(n2061), .Y(n1769) );
    znr3b U896 ( .A(DW6[0]), .B(n2077), .C(n1924), .Y(n1770) );
    znr4b U897 ( .A(UP_DW3[2]), .B(n1839), .C(n2098), .D(n1841), .Y(n1771) );
    znr2b U898 ( .A(n2106), .B(n1991), .Y(n1772) );
    zaoi211b U899 ( .A(n2080), .B(n1931), .C(n1997), .D(n1946), .Y(n1773) );
    zdffqb TCOUNT_reg_0 ( .CK(PCICLK), .D(TCOUNT793_0), .Q(UP_DW5[0]) );
    zivb U900 ( .A(UP_DW5[0]), .Y(n1945) );
    zdffqb RETRYCNT_reg_0 ( .CK(PCICLK), .D(RETRYCNT1095_0), .Q(RETRYCNT_0) );
    zivb U901 ( .A(RETRYCNT_0), .Y(n2119) );
    zor2b U902 ( .A(n1817), .B(UP_DW3[22]), .Y(n1774) );
    ziv11b U903 ( .A(SIDWOFFSET[2]), .Y(n1775), .Z(SIDWOFFSET[1]) );
    ziv11b U904 ( .A(n2176), .Y(TRAN_CMD[8]), .Z(TRAN_CMD[1]) );
    zao211d U905 ( .A(SIDWNUM[2]), .B(PCIEND), .C(SITDSM[3]), .D(n1912), .Y(
        n2166) );
    zan2b U906 ( .A(SITDSM[0]), .B(SITD_PARSE_GO), .Y(n1912) );
    zivc U907 ( .A(n1861), .Y(n1851) );
    zan2b U908 ( .A(n1763), .B(PCIEND), .Y(SITDSMNXT_2) );
    zoa22b U909 ( .A(n1771), .B(n1956), .C(PCIEND), .D(n1957), .Y(n1955) );
    zao21b U910 ( .A(SIDWNUM[2]), .B(PCIEND), .C(n1844), .Y(PARSESITDEND_PRE)
         );
    zivb U911 ( .A(PCIEND), .Y(n1830) );
    zan3b U912 ( .A(n1954), .B(n1964), .C(PCIEND), .Y(n1824) );
    zor2b U913 ( .A(DWCNT[0]), .B(n2168), .Y(n2118) );
    zor3d U914 ( .A(DWCNT[3]), .B(DWCNT[2]), .C(DWCNT[1]), .Y(n2168) );
    zao22b U915 ( .A(UP_DW4[5]), .B(n2170), .C(UP_DW5[5]), .D(n1894), .Y(
        SIHCIADD[5]) );
    zor3d U916 ( .A(DWCNT[3]), .B(DWCNT[2]), .C(DWCNT[1]), .Y(n1894) );
    zivb U917 ( .A(n1832), .Y(n1779) );
    zor2b U918 ( .A(n1779), .B(n1968), .Y(n1901) );
    zor2b U919 ( .A(GEN_PERR), .B(n1955), .Y(n1969) );
    zor2b U920 ( .A(GEN_PERR), .B(n1952), .Y(n1858) );
    zor2b U921 ( .A(GEN_PERR), .B(n1935), .Y(n2085) );
    zivb U922 ( .A(GEN_PERR), .Y(n1832) );
    zor2b U923 ( .A(n2169), .B(n2116), .Y(n2117) );
    zor3d U924 ( .A(DWCNT[3]), .B(DWCNT[2]), .C(DWCNT[1]), .Y(n2169) );
    zivb U925 ( .A(TRAN_CMD[8]), .Y(TRAN_CMD[9]) );
    zor2b U926 ( .A(TRAN_CMD[9]), .B(UP_DW3[1]), .Y(TRAN_CMD[104]) );
    zan2b U927 ( .A(ACTLEN[10]), .B(TRAN_CMD[9]), .Y(_cell_952_U2_Z_10) );
    zoa21b U928 ( .A(TRAN_CMD[9]), .B(n1849), .C(n1851), .Y(n1939) );
    zan3b U929 ( .A(TRAN_CMD[9]), .B(n1983), .C(n1851), .Y(n1982) );
    zmux21hb U930 ( .A(n1748), .B(ACTLEN[9]), .S(n2176), .Y(_cell_952_U2_Z_9)
         );
    zmux21hb U931 ( .A(n1749), .B(ACTLEN[8]), .S(n2176), .Y(_cell_952_U2_Z_8)
         );
    zmux21hb U932 ( .A(n1863), .B(ACTLEN[7]), .S(n2176), .Y(_cell_952_U2_Z_7)
         );
    zmux21hb U933 ( .A(n1747), .B(ACTLEN[6]), .S(n2176), .Y(_cell_952_U2_Z_6)
         );
    zmux21hb U934 ( .A(n1864), .B(ACTLEN[5]), .S(n2176), .Y(_cell_952_U2_Z_5)
         );
    zmux21hb U935 ( .A(n1865), .B(ACTLEN[4]), .S(n2176), .Y(_cell_952_U2_Z_4)
         );
    zmux21hb U936 ( .A(n1866), .B(ACTLEN[3]), .S(n2176), .Y(_cell_952_U2_Z_3)
         );
    zmux21hb U937 ( .A(n1867), .B(ACTLEN[2]), .S(n2176), .Y(_cell_952_U2_Z_2)
         );
    zmux21hb U938 ( .A(n1750), .B(ACTLEN[1]), .S(n2176), .Y(_cell_952_U2_Z_1)
         );
    zmux21hb U939 ( .A(n1746), .B(ACTLEN[0]), .S(n2176), .Y(_cell_952_U2_Z_0)
         );
    zao21b U940 ( .A(n1853), .B(n2176), .C(n1884), .Y(SPLITXSTATE861) );
    zbfd U941 ( .A(UP_DW3[30]), .Y(n1781) );
    zmux21lb U942 ( .A(n2018), .B(n2017), .S(UP_DW3[30]), .Y(TRAN_CMD[91]) );
    zmux21lb U943 ( .A(n2016), .B(n2015), .S(n1781), .Y(TRAN_CMD[92]) );
    zmux21lb U944 ( .A(n2020), .B(n2019), .S(UP_DW3[30]), .Y(TRAN_CMD[90]) );
    zmux21lb U945 ( .A(n2004), .B(n2003), .S(n1781), .Y(TRAN_CMD[98]) );
    zmux21lb U946 ( .A(n2008), .B(n2007), .S(UP_DW3[30]), .Y(TRAN_CMD[96]) );
    zmux21lb U947 ( .A(n2022), .B(n2021), .S(n1781), .Y(TRAN_CMD[89]) );
    zmux21lb U948 ( .A(n2012), .B(n2011), .S(n1781), .Y(TRAN_CMD[94]) );
    zmux21lb U949 ( .A(n2024), .B(n2023), .S(n1781), .Y(TRAN_CMD[88]) );
    zmux21lb U950 ( .A(n2002), .B(n2001), .S(n1781), .Y(TRAN_CMD[99]) );
    zmux21lb U951 ( .A(n2045), .B(n2044), .S(UP_DW3[30]), .Y(TRAN_CMD[100]) );
    zmux21lb U952 ( .A(n2026), .B(n2025), .S(n1781), .Y(TRAN_CMD[87]) );
    zmux21lb U953 ( .A(n2043), .B(n2042), .S(n1781), .Y(TRAN_CMD[101]) );
    zmux21lb U954 ( .A(n2014), .B(n2013), .S(n1781), .Y(TRAN_CMD[93]) );
    zmux21lb U955 ( .A(n2041), .B(n2040), .S(UP_DW3[30]), .Y(TRAN_CMD[102]) );
    zmux21lb U956 ( .A(n2010), .B(n2009), .S(n1781), .Y(TRAN_CMD[95]) );
    zmux21lb U957 ( .A(n2039), .B(n2038), .S(n1781), .Y(TRAN_CMD[103]) );
    zmux21lb U958 ( .A(n2006), .B(n2005), .S(n1781), .Y(TRAN_CMD[97]) );
    zmux21lb U959 ( .A(n2032), .B(n2031), .S(UP_DW3[30]), .Y(TRAN_CMD[84]) );
    zmux21lb U960 ( .A(n2030), .B(n2029), .S(n1781), .Y(TRAN_CMD[85]) );
    zmux21lb U961 ( .A(n2028), .B(n2027), .S(n1781), .Y(TRAN_CMD[86]) );
    zmux21lb U962 ( .A(NDW3_30), .B(UP_DW3[30]), .S(n1851), .Y(n1871) );
    zdffqb PG_reg ( .CK(PCICLK), .D(PG747), .Q(UP_DW3[30]) );
    zao211d U963 ( .A(SIDWNUM[2]), .B(PCIEND), .C(SITDSM[3]), .D(n1912), .Y(
        n1861) );
    zbfd U964 ( .A(n1613), .Y(n1782) );
    zbfd U965 ( .A(n1613), .Y(n1784) );
    zbfb U966 ( .A(n1613), .Y(n1783) );
    zoa211b U967 ( .A(n1857), .B(n1783), .C(n1858), .D(n1837), .Y(BACKSTATE526
        ) );
    zivb U968 ( .A(n1782), .Y(n1838) );
    zdffqrb BACKSTATE_reg ( .CK(PCICLK), .D(BACKSTATE526), .R(TRST_), .Q(n1613
        ) );
    zivb U969 ( .A(TRAN_CMD[8]), .Y(TRAN_CMD[3]) );
    zbfb U970 ( .A(SITDSM[13]), .Y(SIHCIMWR) );
    zdffqrb SITDSM_reg_13 ( .CK(PCICLK), .D(SITDSMNXT_13), .R(TRST_), .Q(
        SITDSM[13]) );
    zivb U971 ( .A(n1775), .Y(SIDWOFFSET[0]) );
    zbfb U972 ( .A(SIDWNUM[2]), .Y(SITDSM[1]) );
    zbfb U973 ( .A(UP_LDW3), .Y(UP_LDW4) );
    zdffqrb_ UP_CACHE_reg ( .CK(PCICLK), .D(UP_CACHE1324), .R(TRST_), .Q(
        UP_LDW3) );
    zbfb U974 ( .A(UP_DW5[12]), .Y(TRAN_CMD[52]) );
    zbfb U975 ( .A(UP_DW5[13]), .Y(TRAN_CMD[53]) );
    zbfb U976 ( .A(UP_DW5[14]), .Y(TRAN_CMD[54]) );
    zbfb U977 ( .A(UP_DW5[15]), .Y(TRAN_CMD[55]) );
    zbfb U978 ( .A(UP_DW5[16]), .Y(TRAN_CMD[56]) );
    zbfb U979 ( .A(UP_DW5[17]), .Y(TRAN_CMD[57]) );
    zbfb U980 ( .A(UP_DW5[18]), .Y(TRAN_CMD[58]) );
    zbfb U981 ( .A(UP_DW5[19]), .Y(TRAN_CMD[59]) );
    zbfb U982 ( .A(UP_DW5[20]), .Y(TRAN_CMD[60]) );
    zbfb U983 ( .A(UP_DW5[21]), .Y(TRAN_CMD[61]) );
    zbfb U984 ( .A(UP_DW5[22]), .Y(TRAN_CMD[62]) );
    zbfb U985 ( .A(UP_DW5[23]), .Y(TRAN_CMD[63]) );
    zbfb U986 ( .A(UP_DW5[24]), .Y(TRAN_CMD[64]) );
    zbfb U987 ( .A(UP_DW5[25]), .Y(TRAN_CMD[65]) );
    zbfb U988 ( .A(UP_DW5[26]), .Y(TRAN_CMD[66]) );
    zbfb U989 ( .A(UP_DW5[27]), .Y(TRAN_CMD[67]) );
    zbfb U990 ( .A(UP_DW5[28]), .Y(TRAN_CMD[68]) );
    zbfb U991 ( .A(UP_DW5[29]), .Y(TRAN_CMD[69]) );
    zbfb U992 ( .A(UP_DW5[30]), .Y(TRAN_CMD[70]) );
    zbfb U993 ( .A(UP_DW5[31]), .Y(TRAN_CMD[71]) );
    zbfb U994 ( .A(UP_DW3[1]), .Y(TRAN_CMD[14]) );
    zbfb U995 ( .A(SIRXERR), .Y(UP_DW3[3]) );
    zdffqrb_ SIRXERR_CUR_reg ( .CK(PCICLK), .D(SIRXERR_CUR1009), .R(TRST_), 
        .Q(SIRXERR) );
    zbfb U996 ( .A(SITDSM[12]), .Y(CACHEPHASE) );
    zdffqrb SITDSM_reg_12 ( .CK(PCICLK), .D(SITDSMNXT_12), .R(TRST_), .Q(
        SITDSM[12]) );
    zbfb U997 ( .A(SITDSM[0]), .Y(SITDIDLE) );
    zdffqsb SITDSM_reg_0 ( .CK(PCICLK), .D(PHASENXT_idle), .S(TRST_), .Q(
        SITDSM[0]) );
    zxo2b U998 ( .A(r203_carry_12), .B(OVERWBOFFSET_12), .Y(
        OVERWBOFFSET_P1150_12) );
    zan2b U999 ( .A(UP_DW4[11]), .B(r203_carry_11), .Y(r203_carry_12) );
    zxo2b U1000 ( .A(UP_DW4[11]), .B(r203_carry_11), .Y(OVERWBOFFSET_P1150_11)
         );
    zan2b U1001 ( .A(_cell_952_U2_Z_0), .B(UP_DW4[0]), .Y(r203_carry_1) );
    zxo2b U1002 ( .A(_cell_952_U2_Z_0), .B(UP_DW4[0]), .Y(OVERWBOFFSET_P1150_0
        ) );
    zxo2b U1003 ( .A(sub_342_carry_10), .B(sub_342_B_not_10), .Y(UNDERFLOW) );
    zor2b U1004 ( .A(UP_DW3[16]), .B(sub_342_B_not_0), .Y(sub_342_carry_1) );
    zxn2b U1005 ( .A(UP_DW3[16]), .B(sub_342_B_not_0), .Y(VIR_TOTALBYTES_0) );
    zymx24hb U1006 ( .A1(DW5[3]), .A2(DW5[2]), .A3(DW5[1]), .A4(DW5[0]), .B1(
        DW12[3]), .B2(DW12[2]), .B3(DW12[1]), .B4(DW12[0]), .S(n1782), .Y1(
        NDW5_3), .Y2(NDW5_2), .Y3(NDW5_1), .Y4(NDW5_0) );
    zymx24hb U1007 ( .A1(DW5[7]), .A2(DW5[6]), .A3(DW5[5]), .A4(DW5[4]), .B1(
        DW12[7]), .B2(DW12[6]), .B3(DW12[5]), .B4(DW12[4]), .S(n1784), .Y1(
        UP_DW5[7]), .Y2(UP_DW5[6]), .Y3(UP_DW5[5]), .Y4(NDW5_4) );
    zymx24hb U1008 ( .A1(DW5[11]), .A2(DW5[10]), .A3(DW5[9]), .A4(DW5[8]), 
        .B1(DW12[11]), .B2(DW12[10]), .B3(DW12[9]), .B4(DW12[8]), .S(n1782), 
        .Y1(UP_DW5[11]), .Y2(UP_DW5[10]), .Y3(UP_DW5[9]), .Y4(UP_DW5[8]) );
    zymx24hb U1009 ( .A1(DW5[15]), .A2(DW5[14]), .A3(DW5[13]), .A4(DW5[12]), 
        .B1(DW12[15]), .B2(DW12[14]), .B3(DW12[13]), .B4(DW12[12]), .S(n1784), 
        .Y1(UP_DW5[15]), .Y2(UP_DW5[14]), .Y3(UP_DW5[13]), .Y4(UP_DW5[12]) );
    zymx24hb U1010 ( .A1(DW5[19]), .A2(DW5[18]), .A3(DW5[17]), .A4(DW5[16]), 
        .B1(DW12[19]), .B2(DW12[18]), .B3(DW12[17]), .B4(DW12[16]), .S(n1784), 
        .Y1(UP_DW5[19]), .Y2(UP_DW5[18]), .Y3(UP_DW5[17]), .Y4(UP_DW5[16]) );
    zymx24hb U1011 ( .A1(DW5[23]), .A2(DW5[22]), .A3(DW5[21]), .A4(DW5[20]), 
        .B1(DW12[23]), .B2(DW12[22]), .B3(DW12[21]), .B4(DW12[20]), .S(n1784), 
        .Y1(UP_DW5[23]), .Y2(UP_DW5[22]), .Y3(UP_DW5[21]), .Y4(UP_DW5[20]) );
    zymx24hb U1012 ( .A1(DW5[27]), .A2(DW5[26]), .A3(DW5[25]), .A4(DW5[24]), 
        .B1(DW12[27]), .B2(DW12[26]), .B3(DW12[25]), .B4(DW12[24]), .S(n1784), 
        .Y1(UP_DW5[27]), .Y2(UP_DW5[26]), .Y3(UP_DW5[25]), .Y4(UP_DW5[24]) );
    zymx24hb U1013 ( .A1(DW5[31]), .A2(DW5[30]), .A3(DW5[29]), .A4(DW5[28]), 
        .B1(DW12[31]), .B2(DW12[30]), .B3(DW12[29]), .B4(DW12[28]), .S(n1784), 
        .Y1(UP_DW5[31]), .Y2(UP_DW5[30]), .Y3(UP_DW5[29]), .Y4(UP_DW5[28]) );
    zmux21hb U1014 ( .A(DW1[0]), .B(DW8[0]), .S(n1782), .Y(TRAN_CMD[33]) );
    zmux21hb U1015 ( .A(DW1[1]), .B(DW8[1]), .S(n1784), .Y(TRAN_CMD[34]) );
    zymx24hb U1016 ( .A1(DW1[5]), .A2(DW1[4]), .A3(DW1[3]), .A4(DW1[2]), .B1(
        DW8[5]), .B2(DW8[4]), .B3(DW8[3]), .B4(DW8[2]), .S(n1782), .Y1(
        TRAN_CMD[38]), .Y2(TRAN_CMD[37]), .Y3(TRAN_CMD[36]), .Y4(TRAN_CMD[35])
         );
    zymx24hb U1017 ( .A1(DW1[10]), .A2(DW1[9]), .A3(DW1[8]), .A4(DW1[6]), .B1(
        DW8[10]), .B2(DW8[9]), .B3(DW8[8]), .B4(DW8[6]), .S(n1784), .Y1(
        TRAN_CMD[31]), .Y2(TRAN_CMD[30]), .Y3(TRAN_CMD[29]), .Y4(TRAN_CMD[39])
         );
    zymx24hb U1018 ( .A1(DW1[18]), .A2(DW1[17]), .A3(DW1[16]), .A4(DW1[11]), 
        .B1(DW8[18]), .B2(DW8[17]), .B3(DW8[16]), .B4(DW8[11]), .S(n1782), 
        .Y1(TRAN_CMD[24]), .Y2(TRAN_CMD[23]), .Y3(TRAN_CMD[22]), .Y4(TRAN_CMD
        [32]) );
    zymx24hb U1019 ( .A1(DW1[22]), .A2(DW1[21]), .A3(DW1[20]), .A4(DW1[19]), 
        .B1(DW8[22]), .B2(DW8[21]), .B3(DW8[20]), .B4(DW8[19]), .S(n1784), 
        .Y1(TRAN_CMD[28]), .Y2(TRAN_CMD[27]), .Y3(TRAN_CMD[26]), .Y4(TRAN_CMD
        [25]) );
    zymx24hb U1020 ( .A1(DW1[27]), .A2(DW1[26]), .A3(DW1[25]), .A4(DW1[24]), 
        .B1(DW8[27]), .B2(DW8[26]), .B3(DW8[25]), .B4(DW8[24]), .S(n1784), 
        .Y1(TRAN_CMD[18]), .Y2(TRAN_CMD[17]), .Y3(TRAN_CMD[16]), .Y4(TRAN_CMD
        [15]) );
    zymx24hd U1021 ( .A1(DW1[31]), .A2(DW1[30]), .A3(DW1[29]), .A4(DW1[28]), 
        .B1(DW8[31]), .B2(DW8[30]), .B3(DW8[29]), .B4(DW8[28]), .S(n1783), 
        .Y1(n2176), .Y2(TRAN_CMD[21]), .Y3(TRAN_CMD[20]), .Y4(TRAN_CMD[19]) );
    zymx24hb U1022 ( .A1(DW4[3]), .A2(DW4[2]), .A3(DW4[1]), .A4(DW4[0]), .B1(
        DW11[3]), .B2(DW11[2]), .B3(DW11[1]), .B4(DW11[0]), .S(n1784), .Y1(
        TRAN_CMD[75]), .Y2(TRAN_CMD[74]), .Y3(TRAN_CMD[73]), .Y4(TRAN_CMD[72])
         );
    zymx24hb U1023 ( .A1(DW4[7]), .A2(DW4[6]), .A3(DW4[5]), .A4(DW4[4]), .B1(
        DW11[7]), .B2(DW11[6]), .B3(DW11[5]), .B4(DW11[4]), .S(n1782), .Y1(
        TRAN_CMD[79]), .Y2(TRAN_CMD[78]), .Y3(TRAN_CMD[77]), .Y4(TRAN_CMD[76])
         );
    zymx24hb U1024 ( .A1(DW4[11]), .A2(DW4[10]), .A3(DW4[9]), .A4(DW4[8]), 
        .B1(DW11[11]), .B2(DW11[10]), .B3(DW11[9]), .B4(DW11[8]), .S(n1782), 
        .Y1(TRAN_CMD[83]), .Y2(TRAN_CMD[82]), .Y3(TRAN_CMD[81]), .Y4(TRAN_CMD
        [80]) );
    zymx24hb U1025 ( .A1(DW4[15]), .A2(DW4[14]), .A3(DW4[13]), .A4(DW4[12]), 
        .B1(DW11[15]), .B2(DW11[14]), .B3(DW11[13]), .B4(DW11[12]), .S(n1782), 
        .Y1(UP_DW4[15]), .Y2(UP_DW4[14]), .Y3(UP_DW4[13]), .Y4(UP_DW4[12]) );
    zymx24hb U1026 ( .A1(DW4[19]), .A2(DW4[18]), .A3(DW4[17]), .A4(DW4[16]), 
        .B1(DW11[19]), .B2(DW11[18]), .B3(DW11[17]), .B4(DW11[16]), .S(n1782), 
        .Y1(UP_DW4[19]), .Y2(UP_DW4[18]), .Y3(UP_DW4[17]), .Y4(UP_DW4[16]) );
    zymx24hb U1027 ( .A1(DW4[23]), .A2(DW4[22]), .A3(DW4[21]), .A4(DW4[20]), 
        .B1(DW11[23]), .B2(DW11[22]), .B3(DW11[21]), .B4(DW11[20]), .S(n1782), 
        .Y1(UP_DW4[23]), .Y2(UP_DW4[22]), .Y3(UP_DW4[21]), .Y4(UP_DW4[20]) );
    zymx24hb U1028 ( .A1(DW4[27]), .A2(DW4[26]), .A3(DW4[25]), .A4(DW4[24]), 
        .B1(DW11[27]), .B2(DW11[26]), .B3(DW11[25]), .B4(DW11[24]), .S(n1782), 
        .Y1(UP_DW4[27]), .Y2(UP_DW4[26]), .Y3(UP_DW4[25]), .Y4(UP_DW4[24]) );
    zymx24hb U1029 ( .A1(DW4[31]), .A2(DW4[30]), .A3(DW4[29]), .A4(DW4[28]), 
        .B1(DW11[31]), .B2(DW11[30]), .B3(DW11[29]), .B4(DW11[28]), .S(n1782), 
        .Y1(UP_DW4[31]), .Y2(UP_DW4[30]), .Y3(UP_DW4[29]), .Y4(UP_DW4[28]) );
    zymx24hb U1030 ( .A1(DW2[3]), .A2(DW2[2]), .A3(DW2[1]), .A4(DW2[0]), .B1(
        DW9[3]), .B2(DW9[2]), .B3(DW9[1]), .B4(DW9[0]), .S(n1782), .Y1(SMASK_3
        ), .Y2(SMASK_2), .Y3(SMASK_1), .Y4(SMASK_0) );
    zymx24hb U1031 ( .A1(DW2[7]), .A2(DW2[6]), .A3(DW2[5]), .A4(DW2[4]), .B1(
        DW9[7]), .B2(DW9[6]), .B3(DW9[5]), .B4(DW9[4]), .S(n1782), .Y1(SMASK_7
        ), .Y2(SMASK_6), .Y3(SMASK_5), .Y4(SMASK_4) );
    zymx24hb U1032 ( .A1(DW2[11]), .A2(DW2[10]), .A3(DW2[9]), .A4(DW2[8]), 
        .B1(DW9[11]), .B2(DW9[10]), .B3(DW9[9]), .B4(DW9[8]), .S(n1784), .Y1(
        CMASK_3), .Y2(CMASK_2), .Y3(CMASK_1), .Y4(CMASK_0) );
    zymx24hb U1033 ( .A1(DW2[15]), .A2(DW2[14]), .A3(DW2[13]), .A4(DW2[12]), 
        .B1(DW9[15]), .B2(DW9[14]), .B3(DW9[13]), .B4(DW9[12]), .S(n1783), 
        .Y1(CMASK_7), .Y2(CMASK_6), .Y3(CMASK_5), .Y4(CMASK_4) );
    zmux21hb U1034 ( .A(DW3[0]), .B(DW10[0]), .S(n1782), .Y(UP_DW3[0]) );
    zmux21hb U1035 ( .A(DW3[1]), .B(DW10[1]), .S(n1783), .Y(SPLITXSTATE_COM)
         );
    zymx24hb U1036 ( .A1(DW3[7]), .A2(DW3[6]), .A3(DW3[4]), .A4(DW3[2]), .B1(
        DW10[7]), .B2(DW10[6]), .B3(DW10[4]), .B4(DW10[2]), .S(n1784), .Y1(
        ACTIVE_COM), .Y2(NDW3_6), .Y3(NDW3_4), .Y4(NDW3_2) );
    zymx24hb U1037 ( .A1(DW3[11]), .A2(DW3[10]), .A3(DW3[9]), .A4(DW3[8]), 
        .B1(DW10[11]), .B2(DW10[10]), .B3(DW10[9]), .B4(DW10[8]), .S(n1782), 
        .Y1(CPROGMASK_COM_3), .Y2(CPROGMASK_COM_2), .Y3(CPROGMASK_COM_1), .Y4(
        CPROGMASK_COM_0) );
    zymx24hb U1038 ( .A1(DW3[15]), .A2(DW3[14]), .A3(DW3[13]), .A4(DW3[12]), 
        .B1(DW10[15]), .B2(DW10[14]), .B3(DW10[13]), .B4(DW10[12]), .S(n1784), 
        .Y1(CPROGMASK_COM_7), .Y2(CPROGMASK_COM_6), .Y3(CPROGMASK_COM_5), .Y4(
        CPROGMASK_COM_4) );
    zymx24hb U1039 ( .A1(DW3[19]), .A2(DW3[18]), .A3(DW3[17]), .A4(DW3[16]), 
        .B1(DW10[19]), .B2(DW10[18]), .B3(DW10[17]), .B4(DW10[16]), .S(n1782), 
        .Y1(NDW3_19), .Y2(NDW3_18), .Y3(NDW3_17), .Y4(NDW3_16) );
    zymx24hb U1040 ( .A1(DW3[23]), .A2(DW3[22]), .A3(DW3[21]), .A4(DW3[20]), 
        .B1(DW10[23]), .B2(DW10[22]), .B3(DW10[21]), .B4(DW10[20]), .S(n1784), 
        .Y1(NDW3_23), .Y2(NDW3_22), .Y3(NDW3_21), .Y4(NDW3_20) );
    zymx24hb U1041 ( .A1(DW3[27]), .A2(DW3[26]), .A3(DW3[25]), .A4(DW3[24]), 
        .B1(DW10[27]), .B2(DW10[26]), .B3(DW10[25]), .B4(DW10[24]), .S(n1784), 
        .Y1(UP_DW3[27]), .Y2(UP_DW3[26]), .Y3(NDW3_25), .Y4(NDW3_24) );
    zymx24hb U1042 ( .A1(DW3[31]), .A2(DW3[30]), .A3(DW3[29]), .A4(DW3[28]), 
        .B1(DW10[31]), .B2(DW10[30]), .B3(DW10[29]), .B4(DW10[28]), .S(n1784), 
        .Y1(UP_DW3[31]), .Y2(NDW3_30), .Y3(UP_DW3[29]), .Y4(UP_DW3[28]) );
    zdffqd SPLITXSTATE_reg ( .CK(PCICLK), .D(SPLITXSTATE861), .Q(UP_DW3[1]) );
    zdffqrd SITDSM_reg_1 ( .CK(PCICLK), .D(SIDWOFFSET[2]), .R(TRST_), .Q(
        SIDWNUM[2]) );
    zfa1b sub_342_U2_6 ( .A(UP_DW3[22]), .B(sub_342_B_not_6), .CI(
        sub_342_carry_6), .CO(sub_342_carry_7), .S(VIR_TOTALBYTES_6) );
    zfa1b sub_342_U2_8 ( .A(UP_DW3[24]), .B(sub_342_B_not_8), .CI(
        sub_342_carry_8), .CO(sub_342_carry_9), .S(VIR_TOTALBYTES_8) );
    zfa1b sub_342_U2_9 ( .A(UP_DW3[25]), .B(sub_342_B_not_9), .CI(
        sub_342_carry_9), .CO(sub_342_carry_10), .S(VIR_TOTALBYTES_9) );
    zfa1b sub_342_U2_1 ( .A(UP_DW3[17]), .B(sub_342_B_not_1), .CI(
        sub_342_carry_1), .CO(sub_342_carry_2), .S(VIR_TOTALBYTES_1) );
    zfa1b sub_342_U2_7 ( .A(UP_DW3[23]), .B(sub_342_B_not_7), .CI(
        sub_342_carry_7), .CO(sub_342_carry_8), .S(VIR_TOTALBYTES_7) );
    zfa1b sub_342_U2_5 ( .A(UP_DW3[21]), .B(sub_342_B_not_5), .CI(
        sub_342_carry_5), .CO(sub_342_carry_6), .S(VIR_TOTALBYTES_5) );
    zfa1b sub_342_U2_3 ( .A(UP_DW3[19]), .B(sub_342_B_not_3), .CI(
        sub_342_carry_3), .CO(sub_342_carry_4), .S(VIR_TOTALBYTES_3) );
    zfa1b sub_342_U2_2 ( .A(UP_DW3[18]), .B(sub_342_B_not_2), .CI(
        sub_342_carry_2), .CO(sub_342_carry_3), .S(VIR_TOTALBYTES_2) );
    zfa1b sub_342_U2_4 ( .A(UP_DW3[20]), .B(sub_342_B_not_4), .CI(
        sub_342_carry_4), .CO(sub_342_carry_5), .S(VIR_TOTALBYTES_4) );
    zfa1b r203_U1_5 ( .A(UP_DW4[5]), .B(_cell_952_U2_Z_5), .CI(r203_carry_5), 
        .CO(r203_carry_6), .S(OVERWBOFFSET_P1150_5) );
    zfa1b r203_U1_4 ( .A(UP_DW4[4]), .B(_cell_952_U2_Z_4), .CI(r203_carry_4), 
        .CO(r203_carry_5), .S(OVERWBOFFSET_P1150_4) );
    zfa1b r203_U1_3 ( .A(UP_DW4[3]), .B(_cell_952_U2_Z_3), .CI(r203_carry_3), 
        .CO(r203_carry_4), .S(OVERWBOFFSET_P1150_3) );
    zfa1b r203_U1_10 ( .A(UP_DW4[10]), .B(_cell_952_U2_Z_10), .CI(
        r203_carry_10), .CO(r203_carry_11), .S(OVERWBOFFSET_P1150_10) );
    zfa1b r203_U1_9 ( .A(UP_DW4[9]), .B(_cell_952_U2_Z_9), .CI(r203_carry_9), 
        .CO(r203_carry_10), .S(OVERWBOFFSET_P1150_9) );
    zfa1b r203_U1_2 ( .A(UP_DW4[2]), .B(_cell_952_U2_Z_2), .CI(r203_carry_2), 
        .CO(r203_carry_3), .S(OVERWBOFFSET_P1150_2) );
    zfa1b r203_U1_7 ( .A(UP_DW4[7]), .B(_cell_952_U2_Z_7), .CI(r203_carry_7), 
        .CO(r203_carry_8), .S(OVERWBOFFSET_P1150_7) );
    zfa1b r203_U1_8 ( .A(UP_DW4[8]), .B(_cell_952_U2_Z_8), .CI(r203_carry_8), 
        .CO(r203_carry_9), .S(OVERWBOFFSET_P1150_8) );
    zfa1b r203_U1_6 ( .A(UP_DW4[6]), .B(_cell_952_U2_Z_6), .CI(r203_carry_6), 
        .CO(r203_carry_7), .S(OVERWBOFFSET_P1150_6) );
    zfa1b r203_U1_1 ( .A(UP_DW4[1]), .B(_cell_952_U2_Z_1), .CI(r203_carry_1), 
        .CO(r203_carry_2), .S(OVERWBOFFSET_P1150_1) );
    zor6b U1043 ( .A(GEN_PERR), .B(n1824), .C(n1825), .D(n1826), .E(n1827), 
        .F(n1828), .Y(PHASENXT_idle) );
    zor3b U1044 ( .A(SITDSM[8]), .B(SITDSM[9]), .C(n1829), .Y(SICMDSTART_P) );
    zao21d U1045 ( .A(n1763), .B(n1830), .C(n1831), .Y(SIDWOFFSET[2]) );
    zan4b U1046 ( .A(TMOUT), .B(n1835), .C(UP_DW3[1]), .D(n2176), .Y(n1834) );
    zan4b U1047 ( .A(n1838), .B(n1839), .C(SITDSM[13]), .D(PCIEND), .Y(
        CACHE_INVALID452) );
    zao211b U1048 ( .A(n1840), .B(n1841), .C(SITDSM[10]), .D(n1842), .Y(
        SIEOT1441) );
    zoa21d U1049 ( .A(SICMDSTART_EOT), .B(SICMDSTART), .C(n1845), .Y(
        SICMDSTART_EOT1404) );
    zor3b U1050 ( .A(n1753), .B(n1859), .C(DW6[2]), .Y(SIHCIADR[2]) );
    zor3b U1051 ( .A(n1753), .B(n2171), .C(DW6[3]), .Y(SIHCIADR[3]) );
    zao222b U1052 ( .A(NDW5_2), .B(n1861), .C(UP_DW5[2]), .D(n1768), .E(
        TCOUNT797_2), .F(n1767), .Y(TCOUNT793_2) );
    zao222b U1053 ( .A(NDW5_1), .B(n1861), .C(n1768), .D(UP_DW5[1]), .E(
        TCOUNT797_1), .F(n1767), .Y(TCOUNT793_1) );
    zao222b U1054 ( .A(NDW5_0), .B(n1861), .C(UP_DW5[0]), .D(n1768), .E(n1945), 
        .F(n1767), .Y(TCOUNT793_0) );
    zao222b U1055 ( .A(UP_DW3[8]), .B(n1872), .C(CPROGMASK_COM_0), .D(n1861), 
        .E(n1873), .F(n1874), .Y(CPROGMASK875_0) );
    zao222b U1056 ( .A(UP_DW3[9]), .B(n1872), .C(CPROGMASK_COM_1), .D(n2166), 
        .E(n1873), .F(n1875), .Y(CPROGMASK875_1) );
    zao222b U1057 ( .A(CPROGMASK_COM_2), .B(n2166), .C(UP_DW3[10]), .D(n1872), 
        .E(n1873), .F(n1876), .Y(CPROGMASK875_2) );
    zao222b U1058 ( .A(CPROGMASK_COM_3), .B(n1861), .C(UP_DW3[11]), .D(n1872), 
        .E(n1873), .F(n1877), .Y(CPROGMASK875_3) );
    zao222b U1059 ( .A(CPROGMASK_COM_4), .B(n2166), .C(UP_DW3[12]), .D(n1872), 
        .E(n1873), .F(n1878), .Y(CPROGMASK875_4) );
    zao222b U1060 ( .A(CPROGMASK_COM_5), .B(n1861), .C(UP_DW3[13]), .D(n1872), 
        .E(n1873), .F(n1879), .Y(CPROGMASK875_5) );
    zao222b U1061 ( .A(CPROGMASK_COM_6), .B(n1861), .C(UP_DW3[14]), .D(n1872), 
        .E(n1873), .F(n1880), .Y(CPROGMASK875_6) );
    zao222b U1062 ( .A(CPROGMASK_COM_7), .B(n1861), .C(UP_DW3[15]), .D(n1872), 
        .E(n1873), .F(n1881), .Y(CPROGMASK875_7) );
    zao211b U1063 ( .A(SITDSM[13]), .B(n1888), .C(n1779), .D(n1889), .Y(
        SITDERRINT_T1552) );
    zao222b U1064 ( .A(NDW5_3), .B(n2166), .C(UP_DW5[3]), .D(n1890), .E(n1891), 
        .F(n1765), .Y(TP757_0) );
    zao222b U1065 ( .A(NDW5_4), .B(n1861), .C(UP_DW5[4]), .D(n1890), .E(n1765), 
        .F(n1892), .Y(TP757_1) );
    zao222b U1066 ( .A(UP_DW3[0]), .B(n2167), .C(UP_DW5[0]), .D(n1894), .E(
        UP_DW4[0]), .F(n1895), .Y(SIHCIADD[0]) );
    zao222b U1067 ( .A(UP_DW5[1]), .B(n2168), .C(n2167), .D(UP_DW3[1]), .E(
        UP_DW4[1]), .F(n2170), .Y(SIHCIADD[1]) );
    zao222b U1068 ( .A(UP_DW5[2]), .B(n2169), .C(UP_DW3[2]), .D(n1893), .E(
        UP_DW4[2]), .F(n1895), .Y(SIHCIADD[2]) );
    zao222b U1069 ( .A(UP_DW5[3]), .B(n1894), .C(SIRXERR), .D(n2167), .E(
        UP_DW4[3]), .F(n2170), .Y(SIHCIADD[3]) );
    zao222b U1070 ( .A(UP_DW5[4]), .B(n2168), .C(UP_DW3[4]), .D(n1893), .E(
        UP_DW4[4]), .F(n1895), .Y(SIHCIADD[4]) );
    zao222b U1071 ( .A(UP_DW3[6]), .B(n1893), .C(UP_DW5[6]), .D(n2168), .E(
        UP_DW4[6]), .F(n2170), .Y(SIHCIADD[6]) );
    zao222b U1072 ( .A(n2167), .B(UP_DW3[7]), .C(UP_DW5[7]), .D(n2169), .E(
        UP_DW4[7]), .F(n1895), .Y(SIHCIADD[7]) );
    zao222b U1073 ( .A(UP_DW3[8]), .B(n2167), .C(UP_DW5[8]), .D(n1894), .E(
        UP_DW4[8]), .F(n2170), .Y(SIHCIADD[8]) );
    zao222b U1074 ( .A(UP_DW3[9]), .B(n1893), .C(UP_DW5[9]), .D(n2168), .E(
        n1895), .F(UP_DW4[9]), .Y(SIHCIADD[9]) );
    zao222b U1075 ( .A(UP_DW3[10]), .B(n2167), .C(UP_DW5[10]), .D(n2169), .E(
        UP_DW4[10]), .F(n1895), .Y(SIHCIADD[10]) );
    zao222b U1076 ( .A(UP_DW3[11]), .B(n1893), .C(UP_DW5[11]), .D(n1894), .E(
        UP_DW4[11]), .F(n2170), .Y(SIHCIADD[11]) );
    zao222b U1077 ( .A(UP_DW5[12]), .B(n2169), .C(UP_DW3[12]), .D(n2167), .E(
        n2170), .F(UP_DW4[12]), .Y(SIHCIADD[12]) );
    zao222b U1078 ( .A(UP_DW5[13]), .B(n1894), .C(UP_DW3[13]), .D(n1893), .E(
        n1895), .F(UP_DW4[13]), .Y(SIHCIADD[13]) );
    zao222b U1079 ( .A(UP_DW5[14]), .B(n2168), .C(UP_DW3[14]), .D(n2167), .E(
        n2170), .F(UP_DW4[14]), .Y(SIHCIADD[14]) );
    zao222b U1080 ( .A(UP_DW5[15]), .B(n2169), .C(UP_DW3[15]), .D(n1893), .E(
        n1895), .F(UP_DW4[15]), .Y(SIHCIADD[15]) );
    zao222b U1081 ( .A(UP_DW5[16]), .B(n1894), .C(n1893), .D(UP_DW3[16]), .E(
        n2170), .F(UP_DW4[16]), .Y(SIHCIADD[16]) );
    zao222b U1082 ( .A(UP_DW5[17]), .B(n2168), .C(n2167), .D(UP_DW3[17]), .E(
        n1895), .F(UP_DW4[17]), .Y(SIHCIADD[17]) );
    zao222b U1083 ( .A(UP_DW5[18]), .B(n2169), .C(n1893), .D(UP_DW3[18]), .E(
        n2170), .F(UP_DW4[18]), .Y(SIHCIADD[18]) );
    zao222b U1084 ( .A(UP_DW5[19]), .B(n1894), .C(n2167), .D(UP_DW3[19]), .E(
        n1895), .F(UP_DW4[19]), .Y(SIHCIADD[19]) );
    zao222b U1085 ( .A(UP_DW5[20]), .B(n2168), .C(n1893), .D(UP_DW3[20]), .E(
        n2170), .F(UP_DW4[20]), .Y(SIHCIADD[20]) );
    zao222b U1086 ( .A(UP_DW5[21]), .B(n2169), .C(n2167), .D(UP_DW3[21]), .E(
        n1895), .F(UP_DW4[21]), .Y(SIHCIADD[21]) );
    zao222b U1087 ( .A(UP_DW5[22]), .B(n1894), .C(n1893), .D(UP_DW3[22]), .E(
        n2170), .F(UP_DW4[22]), .Y(SIHCIADD[22]) );
    zao222b U1088 ( .A(UP_DW5[23]), .B(n2168), .C(n2167), .D(UP_DW3[23]), .E(
        n1895), .F(UP_DW4[23]), .Y(SIHCIADD[23]) );
    zao222b U1089 ( .A(UP_DW5[24]), .B(n2169), .C(n1893), .D(UP_DW3[24]), .E(
        n2170), .F(UP_DW4[24]), .Y(SIHCIADD[24]) );
    zao222b U1090 ( .A(UP_DW5[25]), .B(n1894), .C(n2167), .D(UP_DW3[25]), .E(
        n1895), .F(UP_DW4[25]), .Y(SIHCIADD[25]) );
    zao222b U1091 ( .A(UP_DW5[26]), .B(n2168), .C(UP_DW3[26]), .D(n2167), .E(
        n2170), .F(UP_DW4[26]), .Y(SIHCIADD[26]) );
    zao222b U1092 ( .A(UP_DW5[27]), .B(n2169), .C(UP_DW3[27]), .D(n1893), .E(
        n1895), .F(UP_DW4[27]), .Y(SIHCIADD[27]) );
    zao222b U1093 ( .A(UP_DW5[28]), .B(n1894), .C(UP_DW3[28]), .D(n2167), .E(
        n2170), .F(UP_DW4[28]), .Y(SIHCIADD[28]) );
    zao222b U1094 ( .A(UP_DW5[29]), .B(n2168), .C(UP_DW3[29]), .D(n1893), .E(
        n1895), .F(UP_DW4[29]), .Y(SIHCIADD[29]) );
    zao222b U1095 ( .A(UP_DW5[30]), .B(n2169), .C(n1893), .D(n1781), .E(n2170), 
        .F(UP_DW4[30]), .Y(SIHCIADD[30]) );
    zao222b U1096 ( .A(UP_DW5[31]), .B(n2169), .C(n2167), .D(UP_DW3[31]), .E(
        n1895), .F(UP_DW4[31]), .Y(SIHCIADD[31]) );
    zan4b U1097 ( .A(n1898), .B(n1868), .C(n1899), .D(n1900), .Y(
        SIRXERR_CUR1009) );
    zao222b U1098 ( .A(n1903), .B(UP_DW4[0]), .C(OVERWBOFFSET_P1150_0), .D(
        n1904), .E(TRAN_CMD[72]), .F(n1905), .Y(OVERWBOFFSET1181_0) );
    zao222b U1099 ( .A(n1903), .B(UP_DW4[1]), .C(OVERWBOFFSET_P1150_1), .D(
        n1904), .E(TRAN_CMD[73]), .F(n1905), .Y(OVERWBOFFSET1181_1) );
    zao222b U1100 ( .A(n1903), .B(UP_DW4[2]), .C(OVERWBOFFSET_P1150_2), .D(
        n1904), .E(TRAN_CMD[74]), .F(n1905), .Y(OVERWBOFFSET1181_2) );
    zao222b U1101 ( .A(n1903), .B(UP_DW4[3]), .C(OVERWBOFFSET_P1150_3), .D(
        n1904), .E(TRAN_CMD[75]), .F(n1905), .Y(OVERWBOFFSET1181_3) );
    zao222b U1102 ( .A(n1903), .B(UP_DW4[4]), .C(OVERWBOFFSET_P1150_4), .D(
        n1904), .E(TRAN_CMD[76]), .F(n1905), .Y(OVERWBOFFSET1181_4) );
    zao222b U1103 ( .A(TRAN_CMD[77]), .B(n1905), .C(n1903), .D(UP_DW4[5]), .E(
        OVERWBOFFSET_P1150_5), .F(n1904), .Y(OVERWBOFFSET1181_5) );
    zao222b U1104 ( .A(TRAN_CMD[78]), .B(n1905), .C(n1903), .D(UP_DW4[6]), .E(
        OVERWBOFFSET_P1150_6), .F(n1904), .Y(OVERWBOFFSET1181_6) );
    zao222b U1105 ( .A(TRAN_CMD[79]), .B(n1905), .C(n1903), .D(UP_DW4[7]), .E(
        OVERWBOFFSET_P1150_7), .F(n1904), .Y(OVERWBOFFSET1181_7) );
    zao222b U1106 ( .A(TRAN_CMD[80]), .B(n1905), .C(n1903), .D(UP_DW4[8]), .E(
        OVERWBOFFSET_P1150_8), .F(n1904), .Y(OVERWBOFFSET1181_8) );
    zao222b U1107 ( .A(TRAN_CMD[81]), .B(n1905), .C(n1903), .D(UP_DW4[9]), .E(
        OVERWBOFFSET_P1150_9), .F(n1904), .Y(OVERWBOFFSET1181_9) );
    zao222b U1108 ( .A(TRAN_CMD[82]), .B(n1905), .C(n1903), .D(UP_DW4[10]), 
        .E(OVERWBOFFSET_P1150_10), .F(n1904), .Y(OVERWBOFFSET1181_10) );
    zao222b U1109 ( .A(TRAN_CMD[83]), .B(n1905), .C(n1903), .D(UP_DW4[11]), 
        .E(OVERWBOFFSET_P1150_11), .F(n1904), .Y(OVERWBOFFSET1181_11) );
    zao222b U1110 ( .A(NDW3_25), .B(n2166), .C(UP_DW3[25]), .D(n1907), .E(
        VIR_TOTALBYTES_9), .F(n1762), .Y(TOTALBYTES621_9) );
    zao222b U1111 ( .A(NDW3_24), .B(n1861), .C(UP_DW3[24]), .D(n1907), .E(
        VIR_TOTALBYTES_8), .F(n1762), .Y(TOTALBYTES621_8) );
    zao222b U1112 ( .A(NDW3_23), .B(n2166), .C(UP_DW3[23]), .D(n1907), .E(
        VIR_TOTALBYTES_7), .F(n1762), .Y(TOTALBYTES621_7) );
    zao222b U1113 ( .A(NDW3_22), .B(n2166), .C(UP_DW3[22]), .D(n1907), .E(
        VIR_TOTALBYTES_6), .F(n1762), .Y(TOTALBYTES621_6) );
    zao222b U1114 ( .A(NDW3_21), .B(n2166), .C(UP_DW3[21]), .D(n1907), .E(
        VIR_TOTALBYTES_5), .F(n1762), .Y(TOTALBYTES621_5) );
    zao222b U1115 ( .A(NDW3_20), .B(n2166), .C(UP_DW3[20]), .D(n1907), .E(
        VIR_TOTALBYTES_4), .F(n1762), .Y(TOTALBYTES621_4) );
    zao222b U1116 ( .A(NDW3_19), .B(n2166), .C(UP_DW3[19]), .D(n1907), .E(
        VIR_TOTALBYTES_3), .F(n1762), .Y(TOTALBYTES621_3) );
    zao222b U1117 ( .A(NDW3_18), .B(n2166), .C(UP_DW3[18]), .D(n1907), .E(
        VIR_TOTALBYTES_2), .F(n1762), .Y(TOTALBYTES621_2) );
    zao222b U1118 ( .A(NDW3_17), .B(n2166), .C(UP_DW3[17]), .D(n1907), .E(
        VIR_TOTALBYTES_1), .F(n1762), .Y(TOTALBYTES621_1) );
    zao222b U1119 ( .A(NDW3_16), .B(n2166), .C(UP_DW3[16]), .D(n1907), .E(
        VIR_TOTALBYTES_0), .F(n1762), .Y(TOTALBYTES621_0) );
    zan4b U1120 ( .A(SITDSM[3]), .B(n1908), .C(n1909), .D(n1832), .Y(
        SITDSMNXT_4) );
    zaoi2x4d U1121 ( .A(CMASK_6), .B(n1914), .C(CMASK_7), .D(n1769), .E(
        CMASK_4), .F(n1915), .G(CMASK_5), .H(n1916), .Y(n1913) );
    zaoi2x4d U1122 ( .A(SMASK_6), .B(n1914), .C(SMASK_7), .D(n1769), .E(
        SMASK_4), .F(n1915), .G(SMASK_5), .H(n1916), .Y(n1917) );
    zoa21d U1123 ( .A(SMASK_0), .B(n1925), .C(n1926), .Y(n1924) );
    zoa21d U1124 ( .A(n1926), .B(n1933), .C(n1754), .Y(n1932) );
    zoa21d U1125 ( .A(n1757), .B(n1755), .C(n1841), .Y(n1934) );
    zoa21d U1126 ( .A(SITDSM[3]), .B(n1965), .C(SITDSM[0]), .Y(n1825) );
    zan4b U1127 ( .A(UP_DW3[31]), .B(SITDSM[13]), .C(n1839), .D(n1969), .Y(
        n1968) );
    zan4b U1128 ( .A(n1966), .B(n1832), .C(n1770), .D(n1971), .Y(n1831) );
    zan4b U1129 ( .A(n1972), .B(n1896), .C(n1973), .D(n1974), .Y(n1846) );
    zan4b U1130 ( .A(n1986), .B(n1987), .C(n1988), .D(n1989), .Y(n1985) );
    zoa21d U1131 ( .A(n1985), .B(UNDERFLOW), .C(n1991), .Y(n1990) );
    zor3b U1132 ( .A(SITDSM[7]), .B(SITDSM[5]), .C(n1840), .Y(n2048) );
    zor3b U1133 ( .A(SITDSM[13]), .B(SITDSM[11]), .C(n2047), .Y(n2049) );
    zor3b U1134 ( .A(SITDSM[0]), .B(SIDWNUM[2]), .C(n2050), .Y(n2051) );
    zor3b U1135 ( .A(SITDSM[0]), .B(SITDSM[3]), .C(n1965), .Y(n2054) );
    zor3b U1136 ( .A(SITDSM[7]), .B(n2049), .C(n2055), .Y(n2056) );
    zor3b U1137 ( .A(SIHCIREQ), .B(n2054), .C(n2048), .Y(n2058) );
    zor2d U1138 ( .A(FRNUM[2]), .B(n2067), .Y(n1925) );
    zor5b U1139 ( .A(SIDWNUM[2]), .B(SITDSM[3]), .C(n1868), .D(n1965), .E(
        n2050), .Y(n2079) );
    zor4b U1140 ( .A(SITDSM[4]), .B(SITDSM[3]), .C(n2080), .D(n2051), .Y(n1928
        ) );
    zor4b U1141 ( .A(IMMEDRETRY), .B(n2176), .C(n1943), .D(n1946), .Y(n2096)
         );
    zor3b U1142 ( .A(SITDSM[10]), .B(SITDSM[11]), .C(n2058), .Y(n2097) );
    zor3b U1143 ( .A(SITDSM[9]), .B(n2000), .C(n2097), .Y(n1956) );
    zor3b U1144 ( .A(n1840), .B(n1963), .C(n2056), .Y(n2099) );
    zor5b U1145 ( .A(SITDSM[11]), .B(n2047), .C(n2048), .D(n2103), .E(n2055), 
        .Y(n1957) );
    zor3b U1146 ( .A(RXDATA0), .B(RXDATA1), .C(RXMDATA), .Y(n1941) );
    zor3b U1147 ( .A(RECOVERYMODE), .B(n1882), .C(n1936), .Y(n1967) );
    zor3b U1148 ( .A(n1994), .B(n1839), .C(n2121), .Y(n2120) );
    zor3b U1149 ( .A(n2147), .B(n2148), .C(n2149), .Y(n2146) );
    zao211b U1150 ( .A(n1759), .B(n1888), .C(n1934), .D(n1932), .Y(n1937) );
    zan4b U1151 ( .A(n1945), .B(n1944), .C(n1892), .D(UP_DW5[1]), .Y(n1891) );
    zao222b U1152 ( .A(n2155), .B(n1845), .C(n2156), .D(n1771), .E(n2154), .F(
        n2157), .Y(n2101) );
    zao222b U1153 ( .A(SIDWNUM[2]), .B(n2054), .C(SITDSM[3]), .D(n1965), .E(
        SITDSM[2]), .F(SITDSM[4]), .Y(n1827) );
    zor3b U1154 ( .A(n1746), .B(n1747), .C(n1748), .Y(n1976) );
    zan4b U1155 ( .A(n2094), .B(n2093), .C(n2089), .D(n2088), .Y(n1987) );
    zan4b U1156 ( .A(n2091), .B(n2092), .C(n2090), .D(n2087), .Y(n1988) );
    zor4b U1157 ( .A(n1882), .B(n2079), .C(RECOVERYMODE), .D(n1770), .Y(n1929)
         );
    zoai21d U1158 ( .A(TRAN_CMD[8]), .B(n1983), .C(TRAN_CMD[104]), .Y(n1862)
         );
    zoai21d U1159 ( .A(n1861), .B(n2086), .C(n2123), .Y(n1907) );
    zor3b U1160 ( .A(n1839), .B(n1838), .C(n1969), .Y(n1836) );
    zor4b U1161 ( .A(n1834), .B(CRCERR), .C(PIDERR), .D(n1772), .Y(n2165) );
    zor2d U1162 ( .A(SIDWOFFSET[2]), .B(n1753), .Y(n1860) );
    zao21d U1163 ( .A(n1981), .B(n1853), .C(n2166), .Y(n1905) );
endmodule


module SLAVECTL ( PCICLK, TRST_, SLAVEMODE, SLAVE_ACT, EHCI_MAC_EOT, GEN_PERR, 
    SLBUI_GO, SLHCIREQ, SLCMDSTART, SLADDR, SLREAD, MDO, DATARDY, TDMAEND, 
    SLMAXLEN, PERIOD_CMD, ASYNC_CMD, SL_PERIOD, CRCERR, PIDERR, SL_DATA_PIDERR, 
    SL_ET_ERR, SL_SE_ERR, SL_ACK_ERR, SLAVE_ERR, SL_PCIERR, SL_ERROFFSET );
output [7:0] SLADDR;
input  [31:0] MDO;
output [7:0] SL_ERROFFSET;
output [10:0] SLMAXLEN;
output [31:0] PERIOD_CMD;
output [31:0] ASYNC_CMD;
input  PCICLK, TRST_, SLAVEMODE, EHCI_MAC_EOT, GEN_PERR, DATARDY, TDMAEND, 
    SL_PERIOD, CRCERR, PIDERR, SL_DATA_PIDERR, SL_ET_ERR, SL_SE_ERR, 
    SL_ACK_ERR;
output SLAVE_ACT, SLBUI_GO, SLHCIREQ, SLCMDSTART, SLREAD, SLAVE_ERR, SL_PCIERR;
    wire ASYNC_CMD_PIPE706_30, ASYNC_CMD_PIPE706_17, ASYNC_CMD_PIPE_14, 
        CUR_ASYNCADDR1138_6, CUR_ASYNCADDR_0, PERIOD_CMD_PIPE_20, 
        ASYNC_CMD_PIPE_0, CUR_PERADDR_6, SPAREO6, SL_PCIERR967, 
        ASYNC_CMD744_13, PERIOD_PIPE554_0, PERADDR_4, PERIOD_CMD630_1, 
        ASYNC_CMD744_5, PERIOD_CMD_PIPE592_22, PERIODCMDEXE856, ASYNCADDR465_3, 
        PERIOD_CMD630_27, CUR_ASYNCADDR1113_6, ASYNC_CMD_PIPE706_4, 
        PERIOD_CMD_PIPE592_4, ASYNC_CMD_PIPE_28, PERIOD_CMD630_12, 
        PERIOD_CMD_PIPE592_17, PERIOD_CMD_PIPE_29, ASYNC_CMD_PIPE_9, 
        PERIOD_CMD_PIPE592_30, ASYNC_CMD744_26, PERIOD_CMD_PIPE_15, 
        PERADDR380_6, PERIOD_CMD630_8, CUR_PERADDR1025_5, PERIOD_CMD_PIPE_5, 
        ASYNC_CMD_PIPE_21, SLAVE_ACT232, ASYNC_CMD_PIPE706_22, 
        PERIOD_CMD_PIPE_2, PERIOD_CMD630_29, ASYNC_CMD_PIPE706_25, 
        ASYNC_CMD_PIPE_26, ASYNC_CMD744_21, CUR_PERADDR1025_2, 
        PERIOD_CMD_PIPE_12, PERADDR380_1, SPAREO0_, PERIOD_CMD_PIPE592_10, 
        ASYNCADDR_0, SPAREO8, CUR_PERADDR1050_0, ASYNC_CMD_PIPE706_19, 
        PERIOD_CMD630_15, ASYNCADDR465_4, CUR_ASYNCADDR1113_1, 
        PERIOD_CMD630_20, PERIOD_CMD_PIPE592_3, ASYNC_CMD_PIPE706_3, PERADDR_3, 
        ASYNC_CMD744_28, PERIOD_CMD_PIPE592_25, ASYNC_CMD744_2, 
        PERIOD_CMD_PIPE592_19, PERIOD_CMD630_6, CUR_PERADDR_1, 
        PERIOD_CMD_PIPE_27, ASYNC_CMD_PIPE_7, ASYNC_CMD744_14, SPAREO1, 
        ASYNC_CMD_PIPE_13, CUR_ASYNCADDR1138_1, ASYNC_CMD_PIPE706_10, 
        PERIOD_PIPE_0, ASYNC_CMD_PIPE706_18, ASYNCADDR449_6, PERIOD_CMD630_14, 
        ASYNCADDR_1, PERIOD_CMD_PIPE592_11, SPAREO9, CUR_PERADDR1050_1, 
        ASYNC_CMD744_20, PERIOD_CMD_PIPE_13, CUR_PERADDR1025_3, PERADDR380_0, 
        PERIOD_CMD_PIPE_3, PERIOD_CMD630_28, ASYNC_CMD_PIPE706_24, 
        ASYNC_CMD_PIPE_27, ASYNC_CMD_PIPE_12, CUR_ASYNCADDR1138_0, 
        ASYNC_CMD_PIPE706_11, PERIOD_PIPE_1, CUR_ASYNCADDR_6, 
        PERIOD_CMD_PIPE592_18, CUR_PERADDR_0, PERIOD_CMD_PIPE_26, 
        ASYNC_CMD_PIPE_6, ASYNC_CMD744_15, SPAREO0, PERADDR364_1, PERADDR_2, 
        ASYNC_CMD744_29, PERIOD_CMD_PIPE592_24, ASYNC_CMD744_3, 
        PERIOD_CMD630_7, ASYNCADDR465_5, PERIOD_CMD630_21, SLAVE_ERR930, 
        PERIOD_CMD_PIPE592_2, ASYNC_CMD_PIPE706_2, ASYNCADDR465_2, 
        PERIOD_CMD630_26, ASYNC_CMD_PIPE706_5, PERIOD_CMD_PIPE592_5, 
        ASYNC_CMD_PIPE_29, PERADDR_5, SLSM_2, SLAVE_GO, PERIOD_CMD630_0, 
        ASYNC_CMD744_4, PERIOD_CMD_PIPE592_23, ASYNC_CMD_PIPE_1, 
        PERIOD_CMD_PIPE_21, PERADDR364_6, SPAREO7, ASYNC_CMD744_12, 
        PERIOD_PIPE554_1, SLREAD782, ASYNC_CMD_PIPE706_31, 
        ASYNC_CMD_PIPE706_16, ASYNC_CMD_PIPE_15, SLSMNXT_1, CUR_ASYNCADDR_1, 
        PERIOD_CMD_PIPE_4, ASYNC_CMD_PIPE_20, ASYNC_CMD_PIPE706_23, 
        ASYNC_CMD744_27, PERIOD_CMD_PIPE_14, PERIOD_CMD630_9, 
        CUR_PERADDR1025_4, ASYNCADDR_6, PERIOD_CMD_PIPE592_16, 
        PERIOD_CMD_PIPE_28, ASYNC_CMD_PIPE_8, SLBUI_GO269, 
        PERIOD_CMD_PIPE592_31, CUR_PERADDR1050_6, ASYNCADDR449_1, 
        PERIOD_CMD630_13, CUR_ASYNCADDR_3, PERIOD_CMD630_18, 
        ASYNC_CMD_PIPE706_14, ASYNC_CMD_PIPE_17, CUR_ASYNCADDR1138_5, 
        ASYNC_CMD_PIPE_30, ASYNC_CMD744_10, PERADDR364_4, SPAREO5, 
        CUR_PERADDR_5, PERIOD_CMD_PIPE_23, ASYNC_CMD_PIPE_3, ASYNC_CMD744_6, 
        PERIOD_CMD_PIPE592_21, PERIOD_CMD630_2, ASYNC_PIPE668_1, 
        ASYNC_CMD_PIPE706_28, ASYNC_CMD_PIPE706_7, PERIOD_CMD_PIPE592_7, 
        ASYNCADDR465_0, PERIOD_CMD630_24, CUR_ASYNCADDR1113_5, ASYNCADDR449_3, 
        PERIOD_CMD630_11, ASYNC_FULL, CUR_PERADDR1050_4, ASYNC_CMD744_19, 
        ASYNCADDR_4, PERIOD_CMD_PIPE592_14, PERIOD_CMD_PIPE_16, 
        CUR_PERADDR1025_6, PERIOD_CMD_PIPE592_28, PERIOD_CMD_PIPE_31, 
        PERADDR380_5, SLSM_0, ASYNC_CMD744_25, ASYNC_PIPE_0, ASYNC_CMD_PIPE_22, 
        ASYNC_CMD_PIPE706_21, PERIOD_CMD_PIPE_6, ASYNC_CMD_PIPE706_26, 
        ASYNC_CMD_PIPE_25, ASYNC_CMD_PIPE706_9, PERIOD_CMD_PIPE592_9, 
        PERIOD_CMD_PIPE_1, ASYNC_CMD744_8, PERADDR380_2, CUR_PERADDR1025_1, 
        PERIOD_CMD_PIPE_11, ASYNC_CMD744_22, CUR_PERADDR1050_3, ASYNCADDR_3, 
        PERIOD_CMD_PIPE592_13, ASYNCADDR449_4, PERIOD_CMD630_16, 
        PERIOD_CMD630_31, ASYNC_CMD_PIPE_19, PERIOD_CMD_PIPE592_0, 
        ASYNC_CMD_PIPE706_0, PERIOD_CMD_PIPE_8, CUR_ASYNCADDR1113_2, 
        PERIOD_CMD630_23, PERIOD_CMD_PIPE_18, PERIOD_CMD630_5, 
        PERIOD_CMD_PIPE592_26, ASYNC_CMD744_1, PERADDR_0, SPAREO2, 
        ASYNC_CMD744_30, PERADDR364_3, ASYNC_CMD_PIPE_4, PERIOD_CMD_PIPE_24, 
        ASYNC_CMD744_17, CUR_PERADDR_2, CUR_ASYNCADDR_4, ASYNC_CMD_PIPE_10, 
        CUR_ASYNCADDR1138_2, ASYNC_CMD_PIPE706_13, ASYNCADDR449_5, 
        PERIOD_CMD630_17, PERIOD_CMD630_30, ASYNC_CMD_PIPE_18, 
        CUR_PERADDR1050_2, ASYNCADDR_2, PERIOD_CMD_PIPE592_12, PERADDR380_3, 
        ASYNC_CMD744_9, PERIOD_CMD_PIPE_10, ASYNC_CMD744_23, 
        ASYNC_CMD_PIPE706_27, ASYNC_CMD_PIPE_24, ASYNC_CMD_PIPE706_8, 
        PERIOD_CMD_PIPE592_8, PERIOD_CMD_PIPE_0, CUR_ASYNCADDR_5, 
        ASYNC_CMD_PIPE_11, CUR_ASYNCADDR1138_3, ASYNC_CMD_PIPE706_12, 
        ASYNC_CMD744_31, SPAREO3, PERADDR364_2, ASYNC_CMD744_16, 
        PERIOD_CMD_PIPE_25, SPAREO1_, ASYNC_CMD_PIPE_5, CUR_PERADDR_3, 
        PERIOD_CMD_PIPE_19, PERIOD_CMD630_4, PERIOD_CMD_PIPE592_27, 
        ASYNC_CMD744_0, PERADDR_1, PERIOD_CMD_PIPE592_1, ASYNC_CMD_PIPE706_1, 
        SLHCIREQ306, PERIOD_CMD_PIPE_9, ASYNCADDR465_6, PERIOD_CMD630_22, 
        CUR_ASYNCADDR1113_3, SLAVE_GO156, ASYNC_CMD_PIPE706_29, 
        ASYNC_CMD_PIPE706_6, PERIOD_CMD_PIPE592_6, PERIOD_CMD630_25, 
        ASYNCADDR465_1, CUR_ASYNCADDR1113_4, ASYNC_CMD744_7, 
        PERIOD_CMD_PIPE592_20, ASYNC_PIPE668_0, PERADDR_6, PERIOD_CMD630_3, 
        SLSM_1, ASYNC_CMD744_11, PERADDR364_5, PERIODCMDEXE, SPAREO4, 
        CUR_PERADDR_4, PERIOD_CMD_PIPE_22, ASYNC_CMD_PIPE_2, CUR_ASYNCADDR_2, 
        PERIOD_CMD630_19, SLSMNXT_2, ASYNC_CMD_PIPE706_15, ASYNC_CMD_PIPE_16, 
        CUR_ASYNCADDR1138_4, ASYNC_CMD_PIPE_31, ASYNC_PIPE_1, 
        ASYNC_CMD_PIPE_23, ASYNC_CMD_PIPE706_20, PERIOD_CMD_PIPE_7, 
        PERIOD_CMD_PIPE_17, PERIOD_CMD_PIPE_30, PERIOD_CMD_PIPE592_29, 
        PERADDR380_4, ASYNC_CMD744_24, CUR_PERADDR1050_5, ASYNC_CMD744_18, 
        PERIOD_CMD_PIPE592_15, ASYNCADDR_5, SLAVE_GO_T, ASYNCADDR449_2, 
        PERIOD_CMD630_10, n1641, n1642, n1643, n1644, n1645, n1646, n1647, 
        n1648, n1649, n1650, n1651, add_172_carry_6, add_172_carry_2, 
        add_172_carry_5, add_172_carry_4, add_172_carry_3, add_185_carry_6, 
        add_185_carry_2, add_185_carry_5, add_185_carry_4, add_185_carry_3, 
        add_353_carry_6, add_353_carry_2, add_353_carry_5, add_353_carry_4, 
        add_353_carry_3, add_367_carry_6, add_367_carry_2, add_367_carry_5, 
        add_367_carry_4, add_367_carry_3, n1652, n1653, n1654, n1655, n1656, 
        n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, 
        n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, 
        n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, 
        n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, 
        n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, 
        n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, 
        n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, 
        n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, 
        n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, 
        n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, 
        n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, 
        n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, 
        n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, 
        n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, 
        n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, 
        n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, 
        n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, 
        n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, 
        n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, 
        n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, 
        n1857, n1860;
    assign SLMAXLEN[10] = 1'b1;
    assign SLMAXLEN[9] = 1'b0;
    assign SLMAXLEN[8] = 1'b0;
    assign SLMAXLEN[7] = 1'b0;
    assign SLMAXLEN[6] = 1'b0;
    assign SLMAXLEN[5] = 1'b0;
    assign SLMAXLEN[4] = 1'b0;
    assign SLMAXLEN[3] = 1'b0;
    assign SLMAXLEN[2] = 1'b0;
    assign SLMAXLEN[1] = 1'b0;
    assign SLMAXLEN[0] = 1'b0;
    zaoi211b SPARE592 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE595 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zoai21b SPARE594 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE593 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zdffrb SPARE591 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE598 ( .A(SPAREO5), .Y(SPAREO6) );
    znr3b SPARE596 ( .A(SPAREO2), .B(ASYNC_FULL), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE597 ( .A(SPAREO4), .Y(SPAREO5) );
    zdffrb SPARE590 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE599 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zor2b U673 ( .A(SLSM_0), .B(n1664), .Y(n1749) );
    zor2b U674 ( .A(n1657), .B(n1715), .Y(n1723) );
    zivb U675 ( .A(EHCI_MAC_EOT), .Y(n1715) );
    zivb U676 ( .A(n1723), .Y(n1849) );
    zor2b U677 ( .A(SL_ERROFFSET[7]), .B(n1689), .Y(n1742) );
    zor2b U678 ( .A(n1693), .B(n1716), .Y(n1741) );
    zor2b U679 ( .A(n1691), .B(PERIODCMDEXE), .Y(n1745) );
    zao33b U680 ( .A(n1721), .B(n1725), .C(n1642), .D(SLSM_1), .E(n1655), .F(
        n1726), .Y(n1724) );
    zor2b U681 ( .A(n1717), .B(n1718), .Y(n1721) );
    zor2b U682 ( .A(n1675), .B(n1719), .Y(n1726) );
    zivb U683 ( .A(n1721), .Y(ASYNC_FULL) );
    zan2b U684 ( .A(n1655), .B(n1684), .Y(n1683) );
    zivb U685 ( .A(TDMAEND), .Y(n1684) );
    zmux21lb U686 ( .A(n1749), .B(n1682), .S(SLSM_2), .Y(n1686) );
    zor2b U687 ( .A(n1678), .B(n1694), .Y(n1693) );
    zan3b U688 ( .A(n1679), .B(n1680), .C(n1681), .Y(n1678) );
    zivb U689 ( .A(n1724), .Y(n1681) );
    zor2b U690 ( .A(SLSM_1), .B(n1654), .Y(n1716) );
    zao22b U691 ( .A(n1648), .B(CUR_ASYNCADDR_0), .C(n1714), .D(n1647), .Y(
        CUR_ASYNCADDR1138_0) );
    zao22b U692 ( .A(n1645), .B(CUR_PERADDR_0), .C(n1713), .D(n1644), .Y(
        CUR_PERADDR1050_0) );
    zao22b U693 ( .A(n1665), .B(ASYNCADDR_0), .C(n1737), .D(n1646), .Y(
        ASYNCADDR465_0) );
    zao22b U694 ( .A(n1673), .B(PERADDR_0), .C(n1736), .D(n1666), .Y(
        PERADDR380_0) );
    zivb U695 ( .A(n1687), .Y(SLSMNXT_2) );
    zor2b U696 ( .A(n1674), .B(n1694), .Y(n1687) );
    zao22b U697 ( .A(n1673), .B(PERADDR_6), .C(PERADDR364_6), .D(n1666), .Y(
        PERADDR380_6) );
    zxo2b U698 ( .A(add_172_carry_6), .B(PERADDR_6), .Y(PERADDR364_6) );
    zao22b U699 ( .A(n1673), .B(PERADDR_5), .C(PERADDR364_5), .D(n1666), .Y(
        PERADDR380_5) );
    zhadrb add_172_U1_1_5 ( .A(PERADDR_5), .B(add_172_carry_5), .CO(
        add_172_carry_6), .S(PERADDR364_5) );
    zao22b U700 ( .A(n1673), .B(PERADDR_4), .C(PERADDR364_4), .D(n1666), .Y(
        PERADDR380_4) );
    zhadrb add_172_U1_1_4 ( .A(PERADDR_4), .B(add_172_carry_4), .CO(
        add_172_carry_5), .S(PERADDR364_4) );
    zao22b U701 ( .A(n1673), .B(PERADDR_3), .C(PERADDR364_3), .D(n1666), .Y(
        PERADDR380_3) );
    zhadrb add_172_U1_1_3 ( .A(PERADDR_3), .B(add_172_carry_3), .CO(
        add_172_carry_4), .S(PERADDR364_3) );
    zao22b U702 ( .A(n1673), .B(PERADDR_2), .C(PERADDR364_2), .D(n1666), .Y(
        PERADDR380_2) );
    zhadrb add_172_U1_1_2 ( .A(PERADDR_2), .B(add_172_carry_2), .CO(
        add_172_carry_3), .S(PERADDR364_2) );
    zao22b U703 ( .A(n1673), .B(PERADDR_1), .C(PERADDR364_1), .D(n1666), .Y(
        PERADDR380_1) );
    zivb U704 ( .A(n1738), .Y(n1673) );
    zor2b U705 ( .A(SLBUI_GO), .B(n1857), .Y(n1738) );
    zhadrb add_172_U1_1_1 ( .A(PERADDR_1), .B(PERADDR_0), .CO(add_172_carry_2), 
        .S(PERADDR364_1) );
    zao22b U706 ( .A(n1665), .B(ASYNCADDR_6), .C(ASYNCADDR449_6), .D(n1646), 
        .Y(ASYNCADDR465_6) );
    zxo2b U707 ( .A(add_185_carry_6), .B(ASYNCADDR_6), .Y(ASYNCADDR449_6) );
    zao22b U708 ( .A(n1665), .B(ASYNCADDR_5), .C(ASYNCADDR449_5), .D(n1646), 
        .Y(ASYNCADDR465_5) );
    zhadrb add_185_U1_1_5 ( .A(ASYNCADDR_5), .B(add_185_carry_5), .CO(
        add_185_carry_6), .S(ASYNCADDR449_5) );
    zao22b U709 ( .A(n1665), .B(ASYNCADDR_4), .C(ASYNCADDR449_4), .D(n1646), 
        .Y(ASYNCADDR465_4) );
    zhadrb add_185_U1_1_4 ( .A(ASYNCADDR_4), .B(add_185_carry_4), .CO(
        add_185_carry_5), .S(ASYNCADDR449_4) );
    zao22b U710 ( .A(n1665), .B(ASYNCADDR_3), .C(ASYNCADDR449_3), .D(n1646), 
        .Y(ASYNCADDR465_3) );
    zhadrb add_185_U1_1_3 ( .A(ASYNCADDR_3), .B(add_185_carry_3), .CO(
        add_185_carry_4), .S(ASYNCADDR449_3) );
    zao22b U711 ( .A(n1665), .B(ASYNCADDR_2), .C(ASYNCADDR449_2), .D(n1646), 
        .Y(ASYNCADDR465_2) );
    zhadrb add_185_U1_1_2 ( .A(ASYNCADDR_2), .B(add_185_carry_2), .CO(
        add_185_carry_3), .S(ASYNCADDR449_2) );
    zao22b U712 ( .A(n1665), .B(ASYNCADDR_1), .C(ASYNCADDR449_1), .D(n1646), 
        .Y(ASYNCADDR465_1) );
    zivb U713 ( .A(n1747), .Y(n1665) );
    zhadrb add_185_U1_1_1 ( .A(ASYNCADDR_1), .B(ASYNCADDR_0), .CO(
        add_185_carry_2), .S(ASYNCADDR449_1) );
    zoai21b U714 ( .A(n1670), .B(n1671), .C(n1672), .Y(PERIOD_PIPE554_1) );
    zivb U715 ( .A(n1672), .Y(n1666) );
    zor2b U716 ( .A(SLBUI_GO), .B(n1740), .Y(n1672) );
    zor2b U717 ( .A(PERIOD_PIPE_0), .B(PERIOD_PIPE_1), .Y(n1667) );
    zan3b U718 ( .A(PERIOD_PIPE_1), .B(n1850), .C(PERIODCMDEXE), .Y(n1668) );
    zivb U719 ( .A(n1670), .Y(n1669) );
    zao21b U720 ( .A(n1661), .B(PERIODCMDEXE), .C(n1738), .Y(n1670) );
    zivb U721 ( .A(n1667), .Y(n1720) );
    zmux21lb U722 ( .A(n1762), .B(n1763), .S(n1739), .Y(PERIOD_CMD_PIPE592_31)
         );
    zmux21lb U723 ( .A(n1770), .B(n1771), .S(n1739), .Y(PERIOD_CMD_PIPE592_28)
         );
    zmux21lb U724 ( .A(n1774), .B(n1775), .S(n1651), .Y(PERIOD_CMD_PIPE592_26)
         );
    zmux21lb U725 ( .A(n1778), .B(n1779), .S(n1739), .Y(PERIOD_CMD_PIPE592_24)
         );
    zmux21lb U726 ( .A(n1782), .B(n1783), .S(n1739), .Y(PERIOD_CMD_PIPE592_22)
         );
    zmux21lb U727 ( .A(n1786), .B(n1787), .S(n1739), .Y(PERIOD_CMD_PIPE592_20)
         );
    zmux21lb U728 ( .A(n1790), .B(n1791), .S(n1739), .Y(PERIOD_CMD_PIPE592_19)
         );
    zmux21lb U729 ( .A(n1794), .B(n1795), .S(n1739), .Y(PERIOD_CMD_PIPE592_17)
         );
    zmux21lb U730 ( .A(n1798), .B(n1799), .S(n1651), .Y(PERIOD_CMD_PIPE592_15)
         );
    zmux21lb U731 ( .A(n1802), .B(n1803), .S(n1651), .Y(PERIOD_CMD_PIPE592_13)
         );
    zmux21lb U732 ( .A(n1806), .B(n1807), .S(n1651), .Y(PERIOD_CMD_PIPE592_11)
         );
    zmux21lb U733 ( .A(n1750), .B(n1751), .S(n1651), .Y(PERIOD_CMD_PIPE592_9)
         );
    zmux21lb U734 ( .A(n1754), .B(n1755), .S(n1739), .Y(PERIOD_CMD_PIPE592_7)
         );
    zmux21lb U735 ( .A(n1758), .B(n1759), .S(n1651), .Y(PERIOD_CMD_PIPE592_5)
         );
    zmux21lb U736 ( .A(n1766), .B(n1767), .S(n1651), .Y(PERIOD_CMD_PIPE592_3)
         );
    zmux21lb U737 ( .A(n1810), .B(n1811), .S(n1651), .Y(PERIOD_CMD_PIPE592_1)
         );
    zivb U738 ( .A(n1740), .Y(n1739) );
    zmux21hb U739 ( .A(PERIOD_CMD_PIPE_31), .B(PERIOD_CMD[31]), .S(n1856), .Y(
        PERIOD_CMD630_31) );
    zmux21hb U740 ( .A(PERIOD_CMD_PIPE_30), .B(PERIOD_CMD[30]), .S(n1814), .Y(
        PERIOD_CMD630_30) );
    zmux21hb U741 ( .A(PERIOD_CMD_PIPE_29), .B(PERIOD_CMD[29]), .S(n1814), .Y(
        PERIOD_CMD630_29) );
    zmux21hb U742 ( .A(PERIOD_CMD_PIPE_28), .B(PERIOD_CMD[28]), .S(n1814), .Y(
        PERIOD_CMD630_28) );
    zmux21hb U743 ( .A(PERIOD_CMD_PIPE_27), .B(PERIOD_CMD[27]), .S(n1856), .Y(
        PERIOD_CMD630_27) );
    zmux21hb U744 ( .A(PERIOD_CMD_PIPE_26), .B(PERIOD_CMD[26]), .S(n1856), .Y(
        PERIOD_CMD630_26) );
    zmux21hb U745 ( .A(PERIOD_CMD_PIPE_25), .B(PERIOD_CMD[25]), .S(n1814), .Y(
        PERIOD_CMD630_25) );
    zmux21hb U746 ( .A(PERIOD_CMD_PIPE_24), .B(PERIOD_CMD[24]), .S(n1856), .Y(
        PERIOD_CMD630_24) );
    zmux21hb U747 ( .A(PERIOD_CMD_PIPE_23), .B(PERIOD_CMD[23]), .S(n1814), .Y(
        PERIOD_CMD630_23) );
    zmux21hb U748 ( .A(PERIOD_CMD_PIPE_22), .B(PERIOD_CMD[22]), .S(n1814), .Y(
        PERIOD_CMD630_22) );
    zmux21hb U749 ( .A(PERIOD_CMD_PIPE_21), .B(PERIOD_CMD[21]), .S(n1856), .Y(
        PERIOD_CMD630_21) );
    zmux21hb U750 ( .A(PERIOD_CMD_PIPE_20), .B(PERIOD_CMD[20]), .S(n1856), .Y(
        PERIOD_CMD630_20) );
    zmux21hb U751 ( .A(PERIOD_CMD_PIPE_19), .B(PERIOD_CMD[19]), .S(n1856), .Y(
        PERIOD_CMD630_19) );
    zmux21hb U752 ( .A(PERIOD_CMD_PIPE_18), .B(PERIOD_CMD[18]), .S(n1814), .Y(
        PERIOD_CMD630_18) );
    zmux21hb U753 ( .A(PERIOD_CMD_PIPE_17), .B(PERIOD_CMD[17]), .S(n1856), .Y(
        PERIOD_CMD630_17) );
    zmux21hb U754 ( .A(PERIOD_CMD_PIPE_16), .B(PERIOD_CMD[16]), .S(n1814), .Y(
        PERIOD_CMD630_16) );
    zmux21hb U755 ( .A(PERIOD_CMD_PIPE_15), .B(PERIOD_CMD[15]), .S(n1856), .Y(
        PERIOD_CMD630_15) );
    zmux21hb U756 ( .A(PERIOD_CMD_PIPE_14), .B(PERIOD_CMD[14]), .S(n1814), .Y(
        PERIOD_CMD630_14) );
    zmux21hb U757 ( .A(PERIOD_CMD_PIPE_13), .B(PERIOD_CMD[13]), .S(n1814), .Y(
        PERIOD_CMD630_13) );
    zmux21hb U758 ( .A(PERIOD_CMD_PIPE_12), .B(PERIOD_CMD[12]), .S(n1856), .Y(
        PERIOD_CMD630_12) );
    zmux21hb U759 ( .A(PERIOD_CMD_PIPE_11), .B(PERIOD_CMD[11]), .S(n1856), .Y(
        PERIOD_CMD630_11) );
    zmux21hb U760 ( .A(PERIOD_CMD_PIPE_10), .B(PERIOD_CMD[10]), .S(n1814), .Y(
        PERIOD_CMD630_10) );
    zmux21hb U761 ( .A(PERIOD_CMD_PIPE_9), .B(PERIOD_CMD[9]), .S(n1856), .Y(
        PERIOD_CMD630_9) );
    zmux21hb U762 ( .A(PERIOD_CMD_PIPE_8), .B(PERIOD_CMD[8]), .S(n1814), .Y(
        PERIOD_CMD630_8) );
    zmux21hb U763 ( .A(PERIOD_CMD_PIPE_7), .B(PERIOD_CMD[7]), .S(n1856), .Y(
        PERIOD_CMD630_7) );
    zmux21hb U764 ( .A(PERIOD_CMD_PIPE_6), .B(PERIOD_CMD[6]), .S(n1814), .Y(
        PERIOD_CMD630_6) );
    zmux21hb U765 ( .A(PERIOD_CMD_PIPE_5), .B(PERIOD_CMD[5]), .S(n1856), .Y(
        PERIOD_CMD630_5) );
    zmux21hb U766 ( .A(PERIOD_CMD_PIPE_4), .B(PERIOD_CMD[4]), .S(n1814), .Y(
        PERIOD_CMD630_4) );
    zmux21hb U767 ( .A(PERIOD_CMD_PIPE_3), .B(PERIOD_CMD[3]), .S(n1856), .Y(
        PERIOD_CMD630_3) );
    zmux21hb U768 ( .A(PERIOD_CMD_PIPE_2), .B(PERIOD_CMD[2]), .S(n1814), .Y(
        PERIOD_CMD630_2) );
    zmux21hb U769 ( .A(PERIOD_CMD_PIPE_1), .B(PERIOD_CMD[1]), .S(n1814), .Y(
        PERIOD_CMD630_1) );
    zmux21hb U770 ( .A(PERIOD_CMD_PIPE_0), .B(PERIOD_CMD[0]), .S(n1856), .Y(
        PERIOD_CMD630_0) );
    zivb U771 ( .A(n1852), .Y(n1856) );
    zivb U772 ( .A(n1852), .Y(n1814) );
    zao21b U773 ( .A(n1643), .B(ASYNC_PIPE_1), .C(n1646), .Y(ASYNC_PIPE668_1)
         );
    zor2b U774 ( .A(ASYNC_PIPE_0), .B(ASYNC_PIPE_1), .Y(n1659) );
    zan3b U775 ( .A(n1850), .B(ASYNC_PIPE_1), .C(SL_ERROFFSET[7]), .Y(n1660)
         );
    zor2b U776 ( .A(n1716), .B(n1723), .Y(n1680) );
    zivb U777 ( .A(n1659), .Y(n1675) );
    zivb U778 ( .A(MDO[31]), .Y(n1763) );
    zmux21lb U779 ( .A(n1822), .B(n1765), .S(n1650), .Y(ASYNC_CMD_PIPE706_30)
         );
    zivb U780 ( .A(MDO[30]), .Y(n1765) );
    zmux21lb U781 ( .A(n1824), .B(n1769), .S(n1650), .Y(ASYNC_CMD_PIPE706_29)
         );
    zivb U782 ( .A(MDO[29]), .Y(n1769) );
    zivb U783 ( .A(MDO[28]), .Y(n1771) );
    zmux21lb U784 ( .A(n1826), .B(n1773), .S(n1650), .Y(ASYNC_CMD_PIPE706_27)
         );
    zivb U785 ( .A(MDO[27]), .Y(n1773) );
    zivb U786 ( .A(MDO[26]), .Y(n1775) );
    zmux21lb U787 ( .A(n1828), .B(n1777), .S(n1650), .Y(ASYNC_CMD_PIPE706_25)
         );
    zivb U788 ( .A(MDO[25]), .Y(n1777) );
    zivb U789 ( .A(MDO[24]), .Y(n1779) );
    zmux21lb U790 ( .A(n1830), .B(n1781), .S(n1650), .Y(ASYNC_CMD_PIPE706_23)
         );
    zivb U791 ( .A(MDO[23]), .Y(n1781) );
    zivb U792 ( .A(MDO[22]), .Y(n1783) );
    zmux21lb U793 ( .A(n1832), .B(n1785), .S(n1855), .Y(ASYNC_CMD_PIPE706_21)
         );
    zivb U794 ( .A(MDO[21]), .Y(n1785) );
    zivb U795 ( .A(MDO[20]), .Y(n1787) );
    zivb U796 ( .A(MDO[19]), .Y(n1791) );
    zmux21lb U797 ( .A(n1836), .B(n1793), .S(n1855), .Y(ASYNC_CMD_PIPE706_18)
         );
    zivb U798 ( .A(MDO[18]), .Y(n1793) );
    zivb U799 ( .A(MDO[17]), .Y(n1795) );
    zmux21lb U800 ( .A(n1838), .B(n1797), .S(n1650), .Y(ASYNC_CMD_PIPE706_16)
         );
    zivb U801 ( .A(MDO[16]), .Y(n1797) );
    zivb U802 ( .A(MDO[15]), .Y(n1799) );
    zmux21lb U803 ( .A(n1840), .B(n1801), .S(n1855), .Y(ASYNC_CMD_PIPE706_14)
         );
    zivb U804 ( .A(MDO[14]), .Y(n1801) );
    zivb U805 ( .A(MDO[13]), .Y(n1803) );
    zmux21lb U806 ( .A(n1842), .B(n1805), .S(n1650), .Y(ASYNC_CMD_PIPE706_12)
         );
    zivb U807 ( .A(MDO[12]), .Y(n1805) );
    zivb U808 ( .A(MDO[11]), .Y(n1807) );
    zmux21lb U809 ( .A(n1844), .B(n1809), .S(n1855), .Y(ASYNC_CMD_PIPE706_10)
         );
    zivb U810 ( .A(MDO[10]), .Y(n1809) );
    zivb U811 ( .A(MDO[9]), .Y(n1751) );
    zmux21lb U812 ( .A(n1816), .B(n1753), .S(n1855), .Y(ASYNC_CMD_PIPE706_8)
         );
    zivb U813 ( .A(MDO[8]), .Y(n1753) );
    zivb U814 ( .A(MDO[7]), .Y(n1755) );
    zmux21lb U815 ( .A(n1818), .B(n1757), .S(n1855), .Y(ASYNC_CMD_PIPE706_6)
         );
    zivb U816 ( .A(MDO[6]), .Y(n1757) );
    zivb U817 ( .A(MDO[5]), .Y(n1759) );
    zmux21lb U818 ( .A(n1820), .B(n1761), .S(n1855), .Y(ASYNC_CMD_PIPE706_4)
         );
    zivb U819 ( .A(MDO[4]), .Y(n1761) );
    zivb U820 ( .A(MDO[3]), .Y(n1767) );
    zmux21lb U821 ( .A(n1834), .B(n1789), .S(n1650), .Y(ASYNC_CMD_PIPE706_2)
         );
    zivb U822 ( .A(MDO[2]), .Y(n1789) );
    zivb U823 ( .A(MDO[1]), .Y(n1811) );
    zmux21lb U824 ( .A(n1846), .B(n1813), .S(n1855), .Y(ASYNC_CMD_PIPE706_0)
         );
    zivb U825 ( .A(MDO[0]), .Y(n1813) );
    zivb U826 ( .A(n1676), .Y(n1855) );
    zivb U827 ( .A(DATARDY), .Y(n1719) );
    zmux21hb U828 ( .A(ASYNC_CMD_PIPE_31), .B(ASYNC_CMD[31]), .S(n1854), .Y(
        ASYNC_CMD744_31) );
    zmux21hb U829 ( .A(ASYNC_CMD_PIPE_30), .B(ASYNC_CMD[30]), .S(n1847), .Y(
        ASYNC_CMD744_30) );
    zmux21hb U830 ( .A(ASYNC_CMD_PIPE_29), .B(ASYNC_CMD[29]), .S(n1847), .Y(
        ASYNC_CMD744_29) );
    zmux21hb U831 ( .A(ASYNC_CMD_PIPE_28), .B(ASYNC_CMD[28]), .S(n1847), .Y(
        ASYNC_CMD744_28) );
    zmux21hb U832 ( .A(ASYNC_CMD_PIPE_27), .B(ASYNC_CMD[27]), .S(n1854), .Y(
        ASYNC_CMD744_27) );
    zmux21hb U833 ( .A(ASYNC_CMD_PIPE_26), .B(ASYNC_CMD[26]), .S(n1854), .Y(
        ASYNC_CMD744_26) );
    zmux21hb U834 ( .A(ASYNC_CMD_PIPE_25), .B(ASYNC_CMD[25]), .S(n1847), .Y(
        ASYNC_CMD744_25) );
    zmux21hb U835 ( .A(ASYNC_CMD_PIPE_24), .B(ASYNC_CMD[24]), .S(n1854), .Y(
        ASYNC_CMD744_24) );
    zmux21hb U836 ( .A(ASYNC_CMD_PIPE_23), .B(ASYNC_CMD[23]), .S(n1847), .Y(
        ASYNC_CMD744_23) );
    zmux21hb U837 ( .A(ASYNC_CMD_PIPE_22), .B(ASYNC_CMD[22]), .S(n1847), .Y(
        ASYNC_CMD744_22) );
    zmux21hb U838 ( .A(ASYNC_CMD_PIPE_21), .B(ASYNC_CMD[21]), .S(n1854), .Y(
        ASYNC_CMD744_21) );
    zmux21hb U839 ( .A(ASYNC_CMD_PIPE_20), .B(ASYNC_CMD[20]), .S(n1854), .Y(
        ASYNC_CMD744_20) );
    zmux21hb U840 ( .A(ASYNC_CMD_PIPE_19), .B(ASYNC_CMD[19]), .S(n1854), .Y(
        ASYNC_CMD744_19) );
    zmux21hb U841 ( .A(ASYNC_CMD_PIPE_18), .B(ASYNC_CMD[18]), .S(n1847), .Y(
        ASYNC_CMD744_18) );
    zmux21hb U842 ( .A(ASYNC_CMD_PIPE_17), .B(ASYNC_CMD[17]), .S(n1854), .Y(
        ASYNC_CMD744_17) );
    zmux21hb U843 ( .A(ASYNC_CMD_PIPE_16), .B(ASYNC_CMD[16]), .S(n1847), .Y(
        ASYNC_CMD744_16) );
    zmux21hb U844 ( .A(ASYNC_CMD_PIPE_15), .B(ASYNC_CMD[15]), .S(n1854), .Y(
        ASYNC_CMD744_15) );
    zmux21hb U845 ( .A(ASYNC_CMD_PIPE_14), .B(ASYNC_CMD[14]), .S(n1847), .Y(
        ASYNC_CMD744_14) );
    zmux21hb U846 ( .A(ASYNC_CMD_PIPE_13), .B(ASYNC_CMD[13]), .S(n1847), .Y(
        ASYNC_CMD744_13) );
    zmux21hb U847 ( .A(ASYNC_CMD_PIPE_12), .B(ASYNC_CMD[12]), .S(n1854), .Y(
        ASYNC_CMD744_12) );
    zmux21hb U848 ( .A(ASYNC_CMD_PIPE_11), .B(ASYNC_CMD[11]), .S(n1854), .Y(
        ASYNC_CMD744_11) );
    zmux21hb U849 ( .A(ASYNC_CMD_PIPE_10), .B(ASYNC_CMD[10]), .S(n1847), .Y(
        ASYNC_CMD744_10) );
    zmux21hb U850 ( .A(ASYNC_CMD_PIPE_9), .B(ASYNC_CMD[9]), .S(n1854), .Y(
        ASYNC_CMD744_9) );
    zmux21hb U851 ( .A(ASYNC_CMD_PIPE_8), .B(ASYNC_CMD[8]), .S(n1847), .Y(
        ASYNC_CMD744_8) );
    zmux21hb U852 ( .A(ASYNC_CMD_PIPE_7), .B(ASYNC_CMD[7]), .S(n1854), .Y(
        ASYNC_CMD744_7) );
    zmux21hb U853 ( .A(ASYNC_CMD_PIPE_6), .B(ASYNC_CMD[6]), .S(n1847), .Y(
        ASYNC_CMD744_6) );
    zmux21hb U854 ( .A(ASYNC_CMD_PIPE_5), .B(ASYNC_CMD[5]), .S(n1854), .Y(
        ASYNC_CMD744_5) );
    zmux21hb U855 ( .A(ASYNC_CMD_PIPE_4), .B(ASYNC_CMD[4]), .S(n1847), .Y(
        ASYNC_CMD744_4) );
    zmux21hb U856 ( .A(ASYNC_CMD_PIPE_3), .B(ASYNC_CMD[3]), .S(n1854), .Y(
        ASYNC_CMD744_3) );
    zmux21hb U857 ( .A(ASYNC_CMD_PIPE_2), .B(ASYNC_CMD[2]), .S(n1847), .Y(
        ASYNC_CMD744_2) );
    zmux21hb U858 ( .A(ASYNC_CMD_PIPE_1), .B(ASYNC_CMD[1]), .S(n1847), .Y(
        ASYNC_CMD744_1) );
    zmux21hb U859 ( .A(ASYNC_CMD_PIPE_0), .B(ASYNC_CMD[0]), .S(n1854), .Y(
        ASYNC_CMD744_0) );
    zivb U860 ( .A(n1853), .Y(n1854) );
    zao22b U861 ( .A(n1748), .B(ASYNC_PIPE_1), .C(n1661), .D(SL_ERROFFSET[7]), 
        .Y(n1853) );
    zivb U862 ( .A(n1853), .Y(n1847) );
    zao22b U863 ( .A(n1645), .B(CUR_PERADDR_6), .C(n1644), .D(
        CUR_PERADDR1025_6), .Y(CUR_PERADDR1050_6) );
    zxo2b U864 ( .A(add_353_carry_6), .B(CUR_PERADDR_6), .Y(CUR_PERADDR1025_6)
         );
    zao22b U865 ( .A(n1645), .B(CUR_PERADDR_5), .C(CUR_PERADDR1025_5), .D(
        n1644), .Y(CUR_PERADDR1050_5) );
    zhadrb add_353_U1_1_5 ( .A(CUR_PERADDR_5), .B(add_353_carry_5), .CO(
        add_353_carry_6), .S(CUR_PERADDR1025_5) );
    zao22b U866 ( .A(n1645), .B(CUR_PERADDR_4), .C(CUR_PERADDR1025_4), .D(
        n1644), .Y(CUR_PERADDR1050_4) );
    zhadrb add_353_U1_1_4 ( .A(CUR_PERADDR_4), .B(add_353_carry_4), .CO(
        add_353_carry_5), .S(CUR_PERADDR1025_4) );
    zao22b U867 ( .A(n1645), .B(CUR_PERADDR_3), .C(CUR_PERADDR1025_3), .D(
        n1644), .Y(CUR_PERADDR1050_3) );
    zhadrb add_353_U1_1_3 ( .A(CUR_PERADDR_3), .B(add_353_carry_3), .CO(
        add_353_carry_4), .S(CUR_PERADDR1025_3) );
    zao22b U868 ( .A(n1645), .B(CUR_PERADDR_2), .C(CUR_PERADDR1025_2), .D(
        n1644), .Y(CUR_PERADDR1050_2) );
    zhadrb add_353_U1_1_2 ( .A(CUR_PERADDR_2), .B(add_353_carry_2), .CO(
        add_353_carry_3), .S(CUR_PERADDR1025_2) );
    zao22b U869 ( .A(n1645), .B(CUR_PERADDR_1), .C(CUR_PERADDR1025_1), .D(
        n1644), .Y(CUR_PERADDR1050_1) );
    zivb U870 ( .A(n1742), .Y(n1743) );
    zhadrb add_353_U1_1_1 ( .A(CUR_PERADDR_1), .B(CUR_PERADDR_0), .CO(
        add_353_carry_2), .S(CUR_PERADDR1025_1) );
    zao22b U871 ( .A(n1648), .B(CUR_ASYNCADDR_6), .C(n1647), .D(
        CUR_ASYNCADDR1113_6), .Y(CUR_ASYNCADDR1138_6) );
    zxo2b U872 ( .A(add_367_carry_6), .B(CUR_ASYNCADDR_6), .Y(
        CUR_ASYNCADDR1113_6) );
    zao22b U873 ( .A(n1648), .B(CUR_ASYNCADDR_5), .C(CUR_ASYNCADDR1113_5), .D(
        n1647), .Y(CUR_ASYNCADDR1138_5) );
    zhadrb add_367_U1_1_5 ( .A(CUR_ASYNCADDR_5), .B(add_367_carry_5), .CO(
        add_367_carry_6), .S(CUR_ASYNCADDR1113_5) );
    zao22b U874 ( .A(n1648), .B(CUR_ASYNCADDR_4), .C(CUR_ASYNCADDR1113_4), .D(
        n1647), .Y(CUR_ASYNCADDR1138_4) );
    zhadrb add_367_U1_1_4 ( .A(CUR_ASYNCADDR_4), .B(add_367_carry_4), .CO(
        add_367_carry_5), .S(CUR_ASYNCADDR1113_4) );
    zao22b U875 ( .A(n1648), .B(CUR_ASYNCADDR_3), .C(CUR_ASYNCADDR1113_3), .D(
        n1647), .Y(CUR_ASYNCADDR1138_3) );
    zhadrb add_367_U1_1_3 ( .A(CUR_ASYNCADDR_3), .B(add_367_carry_3), .CO(
        add_367_carry_4), .S(CUR_ASYNCADDR1113_3) );
    zao22b U876 ( .A(n1648), .B(CUR_ASYNCADDR_2), .C(CUR_ASYNCADDR1113_2), .D(
        n1647), .Y(CUR_ASYNCADDR1138_2) );
    zhadrb add_367_U1_1_2 ( .A(CUR_ASYNCADDR_2), .B(add_367_carry_2), .CO(
        add_367_carry_3), .S(CUR_ASYNCADDR1113_2) );
    zao22b U877 ( .A(n1648), .B(CUR_ASYNCADDR_1), .C(CUR_ASYNCADDR1113_1), .D(
        n1647), .Y(CUR_ASYNCADDR1138_1) );
    zivb U878 ( .A(n1745), .Y(n1746) );
    zivb U879 ( .A(n1741), .Y(n1744) );
    zhadrb add_367_U1_1_1 ( .A(CUR_ASYNCADDR_1), .B(CUR_ASYNCADDR_0), .CO(
        add_367_carry_2), .S(CUR_ASYNCADDR1113_1) );
    zivb U880 ( .A(n1694), .Y(n1727) );
    zmux21hb U881 ( .A(PERIODCMDEXE), .B(SL_PERIOD), .S(SLAVE_ACT), .Y(
        PERIODCMDEXE856) );
    zor2b U882 ( .A(n1653), .B(SL_PCIERR), .Y(SL_PCIERR967) );
    zivb U883 ( .A(n1722), .Y(n1655) );
    zor2b U884 ( .A(SLSM_2), .B(n1657), .Y(n1722) );
    zivb U885 ( .A(n1693), .Y(SLSMNXT_1) );
    znr4b U886 ( .A(DATARDY), .B(n1652), .C(SLREAD), .D(SLSM_2), .Y(SLREAD782)
         );
    zan2b U887 ( .A(SLAVE_ACT), .B(n1688), .Y(n1658) );
    zivb U888 ( .A(n1716), .Y(n1851) );
    zcx2b U889 ( .A(SLAVE_GO_T), .B(n1664), .C(n1662), .D(n1663), .Y(
        SLAVE_ERR930) );
    zor2b U890 ( .A(n1703), .B(n1704), .Y(n1662) );
    zivb U891 ( .A(GEN_PERR), .Y(n1703) );
    zivb U892 ( .A(SLAVEMODE), .Y(n1704) );
    zmux21lb U893 ( .A(SLAVE_ERR), .B(n1848), .S(n1661), .Y(n1663) );
    zivb U894 ( .A(n1680), .Y(n1661) );
    zivb U895 ( .A(n1662), .Y(n1653) );
    zmux21lb U896 ( .A(n1714), .B(n1713), .S(PERIODCMDEXE), .Y(SL_ERROFFSET[0]
        ) );
    zmux21lb U897 ( .A(n1702), .B(n1701), .S(PERIODCMDEXE), .Y(SL_ERROFFSET[1]
        ) );
    zmux21lb U898 ( .A(n1712), .B(n1711), .S(PERIODCMDEXE), .Y(SL_ERROFFSET[2]
        ) );
    zmux21lb U899 ( .A(n1710), .B(n1709), .S(PERIODCMDEXE), .Y(SL_ERROFFSET[3]
        ) );
    zmux21lb U900 ( .A(n1700), .B(n1699), .S(PERIODCMDEXE), .Y(SL_ERROFFSET[4]
        ) );
    zmux21lb U901 ( .A(n1708), .B(n1707), .S(PERIODCMDEXE), .Y(SL_ERROFFSET[5]
        ) );
    zmux21lb U902 ( .A(n1706), .B(n1705), .S(PERIODCMDEXE), .Y(SL_ERROFFSET[6]
        ) );
    zmux21lb U903 ( .A(n1737), .B(n1736), .S(n1725), .Y(SLADDR[0]) );
    zmux21lb U904 ( .A(n1698), .B(n1697), .S(n1725), .Y(SLADDR[1]) );
    zmux21lb U905 ( .A(n1735), .B(n1734), .S(n1725), .Y(SLADDR[2]) );
    zmux21lb U906 ( .A(n1733), .B(n1732), .S(n1725), .Y(SLADDR[3]) );
    zmux21lb U907 ( .A(n1696), .B(n1695), .S(n1725), .Y(SLADDR[4]) );
    zmux21lb U908 ( .A(n1731), .B(n1730), .S(n1725), .Y(SLADDR[5]) );
    zmux21lb U909 ( .A(n1729), .B(n1728), .S(n1725), .Y(SLADDR[6]) );
    zivb U910 ( .A(SLADDR[7]), .Y(n1725) );
    zdffqrb SLSM_reg_2 ( .CK(PCICLK), .D(SLSMNXT_2), .R(TRST_), .Q(SLSM_2) );
    zivb U911 ( .A(SLSM_2), .Y(n1654) );
    zdffqrb SLSM_reg_1 ( .CK(PCICLK), .D(SLSMNXT_1), .R(TRST_), .Q(SLSM_1) );
    zivb U912 ( .A(SLSM_1), .Y(n1652) );
    zdffqrb SLSM_reg_0 ( .CK(PCICLK), .D(n1641), .R(TRST_), .Q(SLSM_0) );
    zivb U913 ( .A(SLSM_0), .Y(n1657) );
    zdffqrb PERADDR_reg_6 ( .CK(PCICLK), .D(PERADDR380_6), .R(TRST_), .Q(
        PERADDR_6) );
    zivb U914 ( .A(PERADDR_6), .Y(n1728) );
    zdffqrb PERADDR_reg_5 ( .CK(PCICLK), .D(PERADDR380_5), .R(TRST_), .Q(
        PERADDR_5) );
    zivb U915 ( .A(PERADDR_5), .Y(n1730) );
    zdffqrb PERADDR_reg_4 ( .CK(PCICLK), .D(PERADDR380_4), .R(TRST_), .Q(
        PERADDR_4) );
    zivb U916 ( .A(PERADDR_4), .Y(n1695) );
    zdffqrb PERADDR_reg_3 ( .CK(PCICLK), .D(PERADDR380_3), .R(TRST_), .Q(
        PERADDR_3) );
    zivb U917 ( .A(PERADDR_3), .Y(n1732) );
    zdffqrb PERADDR_reg_2 ( .CK(PCICLK), .D(PERADDR380_2), .R(TRST_), .Q(
        PERADDR_2) );
    zivb U918 ( .A(PERADDR_2), .Y(n1734) );
    zdffqrb PERADDR_reg_1 ( .CK(PCICLK), .D(PERADDR380_1), .R(TRST_), .Q(
        PERADDR_1) );
    zivb U919 ( .A(PERADDR_1), .Y(n1697) );
    zdffqrb ASYNCADDR_reg_6 ( .CK(PCICLK), .D(ASYNCADDR465_6), .R(TRST_), .Q(
        ASYNCADDR_6) );
    zivb U920 ( .A(ASYNCADDR_6), .Y(n1729) );
    zdffqrb ASYNCADDR_reg_5 ( .CK(PCICLK), .D(ASYNCADDR465_5), .R(TRST_), .Q(
        ASYNCADDR_5) );
    zivb U921 ( .A(ASYNCADDR_5), .Y(n1731) );
    zdffqrb ASYNCADDR_reg_4 ( .CK(PCICLK), .D(ASYNCADDR465_4), .R(TRST_), .Q(
        ASYNCADDR_4) );
    zivb U922 ( .A(ASYNCADDR_4), .Y(n1696) );
    zdffqrb ASYNCADDR_reg_3 ( .CK(PCICLK), .D(ASYNCADDR465_3), .R(TRST_), .Q(
        ASYNCADDR_3) );
    zivb U923 ( .A(ASYNCADDR_3), .Y(n1733) );
    zdffqrb ASYNCADDR_reg_2 ( .CK(PCICLK), .D(ASYNCADDR465_2), .R(TRST_), .Q(
        ASYNCADDR_2) );
    zivb U924 ( .A(ASYNCADDR_2), .Y(n1735) );
    zdffqrb ASYNCADDR_reg_1 ( .CK(PCICLK), .D(ASYNCADDR465_1), .R(TRST_), .Q(
        ASYNCADDR_1) );
    zivb U925 ( .A(ASYNCADDR_1), .Y(n1698) );
    zdffrb PERIOD_PIPE_reg_1 ( .CK(PCICLK), .D(PERIOD_PIPE554_1), .R(TRST_), 
        .Q(PERIOD_PIPE_1), .QN(n1671) );
    zdffqrb PERIOD_PIPE_reg_0 ( .CK(PCICLK), .D(PERIOD_PIPE554_0), .R(TRST_), 
        .Q(PERIOD_PIPE_0) );
    zdffqrb PERIOD_CMD_PIPE_reg_31 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_31), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_31) );
    zivb U926 ( .A(PERIOD_CMD_PIPE_31), .Y(n1762) );
    zdffqrb PERIOD_CMD_PIPE_reg_30 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_30), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_30) );
    zivb U927 ( .A(PERIOD_CMD_PIPE_30), .Y(n1764) );
    zdffqrb PERIOD_CMD_PIPE_reg_29 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_29), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_29) );
    zivb U928 ( .A(PERIOD_CMD_PIPE_29), .Y(n1768) );
    zdffqrb PERIOD_CMD_PIPE_reg_28 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_28), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_28) );
    zivb U929 ( .A(PERIOD_CMD_PIPE_28), .Y(n1770) );
    zdffqrb PERIOD_CMD_PIPE_reg_27 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_27), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_27) );
    zivb U930 ( .A(PERIOD_CMD_PIPE_27), .Y(n1772) );
    zdffqrb PERIOD_CMD_PIPE_reg_26 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_26), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_26) );
    zivb U931 ( .A(PERIOD_CMD_PIPE_26), .Y(n1774) );
    zdffqrb PERIOD_CMD_PIPE_reg_25 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_25), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_25) );
    zivb U932 ( .A(PERIOD_CMD_PIPE_25), .Y(n1776) );
    zdffqrb PERIOD_CMD_PIPE_reg_24 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_24), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_24) );
    zivb U933 ( .A(PERIOD_CMD_PIPE_24), .Y(n1778) );
    zdffqrb PERIOD_CMD_PIPE_reg_23 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_23), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_23) );
    zivb U934 ( .A(PERIOD_CMD_PIPE_23), .Y(n1780) );
    zdffqrb PERIOD_CMD_PIPE_reg_22 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_22), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_22) );
    zivb U935 ( .A(PERIOD_CMD_PIPE_22), .Y(n1782) );
    zdffqrb PERIOD_CMD_PIPE_reg_21 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_21), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_21) );
    zivb U936 ( .A(PERIOD_CMD_PIPE_21), .Y(n1784) );
    zdffqrb PERIOD_CMD_PIPE_reg_20 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_20), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_20) );
    zivb U937 ( .A(PERIOD_CMD_PIPE_20), .Y(n1786) );
    zdffqrb PERIOD_CMD_PIPE_reg_19 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_19), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_19) );
    zivb U938 ( .A(PERIOD_CMD_PIPE_19), .Y(n1790) );
    zdffqrb PERIOD_CMD_PIPE_reg_18 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_18), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_18) );
    zivb U939 ( .A(PERIOD_CMD_PIPE_18), .Y(n1792) );
    zdffqrb PERIOD_CMD_PIPE_reg_17 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_17), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_17) );
    zivb U940 ( .A(PERIOD_CMD_PIPE_17), .Y(n1794) );
    zdffqrb PERIOD_CMD_PIPE_reg_16 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_16), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_16) );
    zivb U941 ( .A(PERIOD_CMD_PIPE_16), .Y(n1796) );
    zdffqrb PERIOD_CMD_PIPE_reg_15 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_15), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_15) );
    zivb U942 ( .A(PERIOD_CMD_PIPE_15), .Y(n1798) );
    zdffqrb PERIOD_CMD_PIPE_reg_14 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_14), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_14) );
    zivb U943 ( .A(PERIOD_CMD_PIPE_14), .Y(n1800) );
    zdffqrb PERIOD_CMD_PIPE_reg_13 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_13), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_13) );
    zivb U944 ( .A(PERIOD_CMD_PIPE_13), .Y(n1802) );
    zdffqrb PERIOD_CMD_PIPE_reg_12 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_12), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_12) );
    zivb U945 ( .A(PERIOD_CMD_PIPE_12), .Y(n1804) );
    zdffqrb PERIOD_CMD_PIPE_reg_11 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_11), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_11) );
    zivb U946 ( .A(PERIOD_CMD_PIPE_11), .Y(n1806) );
    zdffqrb PERIOD_CMD_PIPE_reg_10 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_10), 
        .R(TRST_), .Q(PERIOD_CMD_PIPE_10) );
    zivb U947 ( .A(PERIOD_CMD_PIPE_10), .Y(n1808) );
    zdffqrb PERIOD_CMD_PIPE_reg_9 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_9), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_9) );
    zivb U948 ( .A(PERIOD_CMD_PIPE_9), .Y(n1750) );
    zdffqrb PERIOD_CMD_PIPE_reg_8 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_8), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_8) );
    zivb U949 ( .A(PERIOD_CMD_PIPE_8), .Y(n1752) );
    zdffqrb PERIOD_CMD_PIPE_reg_7 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_7), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_7) );
    zivb U950 ( .A(PERIOD_CMD_PIPE_7), .Y(n1754) );
    zdffqrb PERIOD_CMD_PIPE_reg_6 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_6), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_6) );
    zivb U951 ( .A(PERIOD_CMD_PIPE_6), .Y(n1756) );
    zdffqrb PERIOD_CMD_PIPE_reg_5 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_5), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_5) );
    zivb U952 ( .A(PERIOD_CMD_PIPE_5), .Y(n1758) );
    zdffqrb PERIOD_CMD_PIPE_reg_4 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_4), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_4) );
    zivb U953 ( .A(PERIOD_CMD_PIPE_4), .Y(n1760) );
    zdffqrb PERIOD_CMD_PIPE_reg_3 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_3), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_3) );
    zivb U954 ( .A(PERIOD_CMD_PIPE_3), .Y(n1766) );
    zdffqrb PERIOD_CMD_PIPE_reg_2 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_2), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_2) );
    zivb U955 ( .A(PERIOD_CMD_PIPE_2), .Y(n1788) );
    zdffqrb PERIOD_CMD_PIPE_reg_1 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_1), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_1) );
    zivb U956 ( .A(PERIOD_CMD_PIPE_1), .Y(n1810) );
    zdffqrb PERIOD_CMD_PIPE_reg_0 ( .CK(PCICLK), .D(PERIOD_CMD_PIPE592_0), .R(
        TRST_), .Q(PERIOD_CMD_PIPE_0) );
    zivb U957 ( .A(PERIOD_CMD_PIPE_0), .Y(n1812) );
    zdffqrb PERIOD_CMD_reg_31 ( .CK(PCICLK), .D(PERIOD_CMD630_31), .R(TRST_), 
        .Q(PERIOD_CMD[31]) );
    zdffqrb PERIOD_CMD_reg_30 ( .CK(PCICLK), .D(PERIOD_CMD630_30), .R(TRST_), 
        .Q(PERIOD_CMD[30]) );
    zdffqrb PERIOD_CMD_reg_29 ( .CK(PCICLK), .D(PERIOD_CMD630_29), .R(TRST_), 
        .Q(PERIOD_CMD[29]) );
    zdffqrb PERIOD_CMD_reg_28 ( .CK(PCICLK), .D(PERIOD_CMD630_28), .R(TRST_), 
        .Q(PERIOD_CMD[28]) );
    zdffqrb PERIOD_CMD_reg_27 ( .CK(PCICLK), .D(PERIOD_CMD630_27), .R(TRST_), 
        .Q(PERIOD_CMD[27]) );
    zdffqrb PERIOD_CMD_reg_26 ( .CK(PCICLK), .D(PERIOD_CMD630_26), .R(TRST_), 
        .Q(PERIOD_CMD[26]) );
    zdffqrb PERIOD_CMD_reg_25 ( .CK(PCICLK), .D(PERIOD_CMD630_25), .R(TRST_), 
        .Q(PERIOD_CMD[25]) );
    zdffqrb PERIOD_CMD_reg_24 ( .CK(PCICLK), .D(PERIOD_CMD630_24), .R(TRST_), 
        .Q(PERIOD_CMD[24]) );
    zdffqrb PERIOD_CMD_reg_23 ( .CK(PCICLK), .D(PERIOD_CMD630_23), .R(TRST_), 
        .Q(PERIOD_CMD[23]) );
    zdffqrb PERIOD_CMD_reg_22 ( .CK(PCICLK), .D(PERIOD_CMD630_22), .R(TRST_), 
        .Q(PERIOD_CMD[22]) );
    zdffqrb PERIOD_CMD_reg_21 ( .CK(PCICLK), .D(PERIOD_CMD630_21), .R(TRST_), 
        .Q(PERIOD_CMD[21]) );
    zdffqrb PERIOD_CMD_reg_20 ( .CK(PCICLK), .D(PERIOD_CMD630_20), .R(TRST_), 
        .Q(PERIOD_CMD[20]) );
    zdffqrb PERIOD_CMD_reg_19 ( .CK(PCICLK), .D(PERIOD_CMD630_19), .R(TRST_), 
        .Q(PERIOD_CMD[19]) );
    zdffqrb PERIOD_CMD_reg_18 ( .CK(PCICLK), .D(PERIOD_CMD630_18), .R(TRST_), 
        .Q(PERIOD_CMD[18]) );
    zdffqrb PERIOD_CMD_reg_17 ( .CK(PCICLK), .D(PERIOD_CMD630_17), .R(TRST_), 
        .Q(PERIOD_CMD[17]) );
    zdffqrb PERIOD_CMD_reg_16 ( .CK(PCICLK), .D(PERIOD_CMD630_16), .R(TRST_), 
        .Q(PERIOD_CMD[16]) );
    zdffqrb PERIOD_CMD_reg_15 ( .CK(PCICLK), .D(PERIOD_CMD630_15), .R(TRST_), 
        .Q(PERIOD_CMD[15]) );
    zdffqrb PERIOD_CMD_reg_14 ( .CK(PCICLK), .D(PERIOD_CMD630_14), .R(TRST_), 
        .Q(PERIOD_CMD[14]) );
    zdffqrb PERIOD_CMD_reg_13 ( .CK(PCICLK), .D(PERIOD_CMD630_13), .R(TRST_), 
        .Q(PERIOD_CMD[13]) );
    zdffqrb PERIOD_CMD_reg_12 ( .CK(PCICLK), .D(PERIOD_CMD630_12), .R(TRST_), 
        .Q(PERIOD_CMD[12]) );
    zdffqrb PERIOD_CMD_reg_11 ( .CK(PCICLK), .D(PERIOD_CMD630_11), .R(TRST_), 
        .Q(PERIOD_CMD[11]) );
    zdffqrb PERIOD_CMD_reg_10 ( .CK(PCICLK), .D(PERIOD_CMD630_10), .R(TRST_), 
        .Q(PERIOD_CMD[10]) );
    zdffqrb PERIOD_CMD_reg_9 ( .CK(PCICLK), .D(PERIOD_CMD630_9), .R(TRST_), 
        .Q(PERIOD_CMD[9]) );
    zdffqrb PERIOD_CMD_reg_8 ( .CK(PCICLK), .D(PERIOD_CMD630_8), .R(TRST_), 
        .Q(PERIOD_CMD[8]) );
    zdffqrb PERIOD_CMD_reg_7 ( .CK(PCICLK), .D(PERIOD_CMD630_7), .R(TRST_), 
        .Q(PERIOD_CMD[7]) );
    zdffqrb PERIOD_CMD_reg_6 ( .CK(PCICLK), .D(PERIOD_CMD630_6), .R(TRST_), 
        .Q(PERIOD_CMD[6]) );
    zdffqrb PERIOD_CMD_reg_5 ( .CK(PCICLK), .D(PERIOD_CMD630_5), .R(TRST_), 
        .Q(PERIOD_CMD[5]) );
    zdffqrb PERIOD_CMD_reg_4 ( .CK(PCICLK), .D(PERIOD_CMD630_4), .R(TRST_), 
        .Q(PERIOD_CMD[4]) );
    zdffqrb PERIOD_CMD_reg_3 ( .CK(PCICLK), .D(PERIOD_CMD630_3), .R(TRST_), 
        .Q(PERIOD_CMD[3]) );
    zdffqrb PERIOD_CMD_reg_2 ( .CK(PCICLK), .D(PERIOD_CMD630_2), .R(TRST_), 
        .Q(PERIOD_CMD[2]) );
    zdffqrb PERIOD_CMD_reg_1 ( .CK(PCICLK), .D(PERIOD_CMD630_1), .R(TRST_), 
        .Q(PERIOD_CMD[1]) );
    zdffqrb PERIOD_CMD_reg_0 ( .CK(PCICLK), .D(PERIOD_CMD630_0), .R(TRST_), 
        .Q(PERIOD_CMD[0]) );
    zdffqrb ASYNC_PIPE_reg_1 ( .CK(PCICLK), .D(ASYNC_PIPE668_1), .R(TRST_), 
        .Q(ASYNC_PIPE_1) );
    zivb U958 ( .A(ASYNC_PIPE_1), .Y(n1718) );
    zdffqrb ASYNC_PIPE_reg_0 ( .CK(PCICLK), .D(ASYNC_PIPE668_0), .R(TRST_), 
        .Q(ASYNC_PIPE_0) );
    zivb U959 ( .A(ASYNC_PIPE_0), .Y(n1717) );
    zdffqrb ASYNC_CMD_PIPE_reg_31 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_31), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_31) );
    zivb U960 ( .A(ASYNC_CMD_PIPE_31), .Y(n1821) );
    zdffqrb ASYNC_CMD_PIPE_reg_30 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_30), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_30) );
    zivb U961 ( .A(ASYNC_CMD_PIPE_30), .Y(n1822) );
    zdffqrb ASYNC_CMD_PIPE_reg_29 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_29), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_29) );
    zivb U962 ( .A(ASYNC_CMD_PIPE_29), .Y(n1824) );
    zdffqrb ASYNC_CMD_PIPE_reg_28 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_28), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_28) );
    zivb U963 ( .A(ASYNC_CMD_PIPE_28), .Y(n1825) );
    zdffqrb ASYNC_CMD_PIPE_reg_27 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_27), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_27) );
    zivb U964 ( .A(ASYNC_CMD_PIPE_27), .Y(n1826) );
    zdffqrb ASYNC_CMD_PIPE_reg_26 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_26), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_26) );
    zivb U965 ( .A(ASYNC_CMD_PIPE_26), .Y(n1827) );
    zdffqrb ASYNC_CMD_PIPE_reg_25 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_25), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_25) );
    zivb U966 ( .A(ASYNC_CMD_PIPE_25), .Y(n1828) );
    zdffqrb ASYNC_CMD_PIPE_reg_24 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_24), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_24) );
    zivb U967 ( .A(ASYNC_CMD_PIPE_24), .Y(n1829) );
    zdffqrb ASYNC_CMD_PIPE_reg_23 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_23), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_23) );
    zivb U968 ( .A(ASYNC_CMD_PIPE_23), .Y(n1830) );
    zdffqrb ASYNC_CMD_PIPE_reg_22 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_22), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_22) );
    zivb U969 ( .A(ASYNC_CMD_PIPE_22), .Y(n1831) );
    zdffqrb ASYNC_CMD_PIPE_reg_21 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_21), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_21) );
    zivb U970 ( .A(ASYNC_CMD_PIPE_21), .Y(n1832) );
    zdffqrb ASYNC_CMD_PIPE_reg_20 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_20), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_20) );
    zivb U971 ( .A(ASYNC_CMD_PIPE_20), .Y(n1833) );
    zdffqrb ASYNC_CMD_PIPE_reg_19 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_19), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_19) );
    zivb U972 ( .A(ASYNC_CMD_PIPE_19), .Y(n1835) );
    zdffqrb ASYNC_CMD_PIPE_reg_18 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_18), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_18) );
    zivb U973 ( .A(ASYNC_CMD_PIPE_18), .Y(n1836) );
    zdffqrb ASYNC_CMD_PIPE_reg_17 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_17), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_17) );
    zivb U974 ( .A(ASYNC_CMD_PIPE_17), .Y(n1837) );
    zdffqrb ASYNC_CMD_PIPE_reg_16 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_16), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_16) );
    zivb U975 ( .A(ASYNC_CMD_PIPE_16), .Y(n1838) );
    zdffqrb ASYNC_CMD_PIPE_reg_15 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_15), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_15) );
    zivb U976 ( .A(ASYNC_CMD_PIPE_15), .Y(n1839) );
    zdffqrb ASYNC_CMD_PIPE_reg_14 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_14), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_14) );
    zivb U977 ( .A(ASYNC_CMD_PIPE_14), .Y(n1840) );
    zdffqrb ASYNC_CMD_PIPE_reg_13 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_13), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_13) );
    zivb U978 ( .A(ASYNC_CMD_PIPE_13), .Y(n1841) );
    zdffqrb ASYNC_CMD_PIPE_reg_12 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_12), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_12) );
    zivb U979 ( .A(ASYNC_CMD_PIPE_12), .Y(n1842) );
    zdffqrb ASYNC_CMD_PIPE_reg_11 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_11), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_11) );
    zivb U980 ( .A(ASYNC_CMD_PIPE_11), .Y(n1843) );
    zdffqrb ASYNC_CMD_PIPE_reg_10 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_10), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_10) );
    zivb U981 ( .A(ASYNC_CMD_PIPE_10), .Y(n1844) );
    zdffqrb ASYNC_CMD_PIPE_reg_9 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_9), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_9) );
    zivb U982 ( .A(ASYNC_CMD_PIPE_9), .Y(n1815) );
    zdffqrb ASYNC_CMD_PIPE_reg_8 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_8), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_8) );
    zivb U983 ( .A(ASYNC_CMD_PIPE_8), .Y(n1816) );
    zdffqrb ASYNC_CMD_PIPE_reg_7 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_7), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_7) );
    zivb U984 ( .A(ASYNC_CMD_PIPE_7), .Y(n1817) );
    zdffqrb ASYNC_CMD_PIPE_reg_6 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_6), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_6) );
    zivb U985 ( .A(ASYNC_CMD_PIPE_6), .Y(n1818) );
    zdffqrb ASYNC_CMD_PIPE_reg_5 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_5), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_5) );
    zivb U986 ( .A(ASYNC_CMD_PIPE_5), .Y(n1819) );
    zdffqrb ASYNC_CMD_PIPE_reg_4 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_4), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_4) );
    zivb U987 ( .A(ASYNC_CMD_PIPE_4), .Y(n1820) );
    zdffqrb ASYNC_CMD_PIPE_reg_3 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_3), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_3) );
    zivb U988 ( .A(ASYNC_CMD_PIPE_3), .Y(n1823) );
    zdffqrb ASYNC_CMD_PIPE_reg_2 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_2), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_2) );
    zivb U989 ( .A(ASYNC_CMD_PIPE_2), .Y(n1834) );
    zdffqrb ASYNC_CMD_PIPE_reg_1 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_1), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_1) );
    zivb U990 ( .A(ASYNC_CMD_PIPE_1), .Y(n1845) );
    zdffqrb ASYNC_CMD_PIPE_reg_0 ( .CK(PCICLK), .D(ASYNC_CMD_PIPE706_0), .R(
        TRST_), .Q(ASYNC_CMD_PIPE_0) );
    zivb U991 ( .A(ASYNC_CMD_PIPE_0), .Y(n1846) );
    zdffqrb ASYNC_CMD_reg_31 ( .CK(PCICLK), .D(ASYNC_CMD744_31), .R(TRST_), 
        .Q(ASYNC_CMD[31]) );
    zdffqrb ASYNC_CMD_reg_30 ( .CK(PCICLK), .D(ASYNC_CMD744_30), .R(TRST_), 
        .Q(ASYNC_CMD[30]) );
    zdffqrb ASYNC_CMD_reg_29 ( .CK(PCICLK), .D(ASYNC_CMD744_29), .R(TRST_), 
        .Q(ASYNC_CMD[29]) );
    zdffqrb ASYNC_CMD_reg_28 ( .CK(PCICLK), .D(ASYNC_CMD744_28), .R(TRST_), 
        .Q(ASYNC_CMD[28]) );
    zdffqrb ASYNC_CMD_reg_27 ( .CK(PCICLK), .D(ASYNC_CMD744_27), .R(TRST_), 
        .Q(ASYNC_CMD[27]) );
    zdffqrb ASYNC_CMD_reg_26 ( .CK(PCICLK), .D(ASYNC_CMD744_26), .R(TRST_), 
        .Q(ASYNC_CMD[26]) );
    zdffqrb ASYNC_CMD_reg_25 ( .CK(PCICLK), .D(ASYNC_CMD744_25), .R(TRST_), 
        .Q(ASYNC_CMD[25]) );
    zdffqrb ASYNC_CMD_reg_24 ( .CK(PCICLK), .D(ASYNC_CMD744_24), .R(TRST_), 
        .Q(ASYNC_CMD[24]) );
    zdffqrb ASYNC_CMD_reg_23 ( .CK(PCICLK), .D(ASYNC_CMD744_23), .R(TRST_), 
        .Q(ASYNC_CMD[23]) );
    zdffqrb ASYNC_CMD_reg_22 ( .CK(PCICLK), .D(ASYNC_CMD744_22), .R(TRST_), 
        .Q(ASYNC_CMD[22]) );
    zdffqrb ASYNC_CMD_reg_21 ( .CK(PCICLK), .D(ASYNC_CMD744_21), .R(TRST_), 
        .Q(ASYNC_CMD[21]) );
    zdffqrb ASYNC_CMD_reg_20 ( .CK(PCICLK), .D(ASYNC_CMD744_20), .R(TRST_), 
        .Q(ASYNC_CMD[20]) );
    zdffqrb ASYNC_CMD_reg_19 ( .CK(PCICLK), .D(ASYNC_CMD744_19), .R(TRST_), 
        .Q(ASYNC_CMD[19]) );
    zdffqrb ASYNC_CMD_reg_18 ( .CK(PCICLK), .D(ASYNC_CMD744_18), .R(TRST_), 
        .Q(ASYNC_CMD[18]) );
    zdffqrb ASYNC_CMD_reg_17 ( .CK(PCICLK), .D(ASYNC_CMD744_17), .R(TRST_), 
        .Q(ASYNC_CMD[17]) );
    zdffqrb ASYNC_CMD_reg_16 ( .CK(PCICLK), .D(ASYNC_CMD744_16), .R(TRST_), 
        .Q(ASYNC_CMD[16]) );
    zdffqrb ASYNC_CMD_reg_15 ( .CK(PCICLK), .D(ASYNC_CMD744_15), .R(TRST_), 
        .Q(ASYNC_CMD[15]) );
    zdffqrb ASYNC_CMD_reg_14 ( .CK(PCICLK), .D(ASYNC_CMD744_14), .R(TRST_), 
        .Q(ASYNC_CMD[14]) );
    zdffqrb ASYNC_CMD_reg_13 ( .CK(PCICLK), .D(ASYNC_CMD744_13), .R(TRST_), 
        .Q(ASYNC_CMD[13]) );
    zdffqrb ASYNC_CMD_reg_12 ( .CK(PCICLK), .D(ASYNC_CMD744_12), .R(TRST_), 
        .Q(ASYNC_CMD[12]) );
    zdffqrb ASYNC_CMD_reg_11 ( .CK(PCICLK), .D(ASYNC_CMD744_11), .R(TRST_), 
        .Q(ASYNC_CMD[11]) );
    zdffqrb ASYNC_CMD_reg_10 ( .CK(PCICLK), .D(ASYNC_CMD744_10), .R(TRST_), 
        .Q(ASYNC_CMD[10]) );
    zdffqrb ASYNC_CMD_reg_9 ( .CK(PCICLK), .D(ASYNC_CMD744_9), .R(TRST_), .Q(
        ASYNC_CMD[9]) );
    zdffqrb ASYNC_CMD_reg_8 ( .CK(PCICLK), .D(ASYNC_CMD744_8), .R(TRST_), .Q(
        ASYNC_CMD[8]) );
    zdffqrb ASYNC_CMD_reg_7 ( .CK(PCICLK), .D(ASYNC_CMD744_7), .R(TRST_), .Q(
        ASYNC_CMD[7]) );
    zdffqrb ASYNC_CMD_reg_6 ( .CK(PCICLK), .D(ASYNC_CMD744_6), .R(TRST_), .Q(
        ASYNC_CMD[6]) );
    zdffqrb ASYNC_CMD_reg_5 ( .CK(PCICLK), .D(ASYNC_CMD744_5), .R(TRST_), .Q(
        ASYNC_CMD[5]) );
    zdffqrb ASYNC_CMD_reg_4 ( .CK(PCICLK), .D(ASYNC_CMD744_4), .R(TRST_), .Q(
        ASYNC_CMD[4]) );
    zdffqrb ASYNC_CMD_reg_3 ( .CK(PCICLK), .D(ASYNC_CMD744_3), .R(TRST_), .Q(
        ASYNC_CMD[3]) );
    zdffqrb ASYNC_CMD_reg_2 ( .CK(PCICLK), .D(ASYNC_CMD744_2), .R(TRST_), .Q(
        ASYNC_CMD[2]) );
    zdffqrb ASYNC_CMD_reg_1 ( .CK(PCICLK), .D(ASYNC_CMD744_1), .R(TRST_), .Q(
        ASYNC_CMD[1]) );
    zdffqrb ASYNC_CMD_reg_0 ( .CK(PCICLK), .D(ASYNC_CMD744_0), .R(TRST_), .Q(
        ASYNC_CMD[0]) );
    zdffqrb CUR_PERADDR_reg_6 ( .CK(PCICLK), .D(CUR_PERADDR1050_6), .R(TRST_), 
        .Q(CUR_PERADDR_6) );
    zivb U992 ( .A(CUR_PERADDR_6), .Y(n1705) );
    zdffqrb CUR_PERADDR_reg_5 ( .CK(PCICLK), .D(CUR_PERADDR1050_5), .R(TRST_), 
        .Q(CUR_PERADDR_5) );
    zivb U993 ( .A(CUR_PERADDR_5), .Y(n1707) );
    zdffqrb CUR_PERADDR_reg_4 ( .CK(PCICLK), .D(CUR_PERADDR1050_4), .R(TRST_), 
        .Q(CUR_PERADDR_4) );
    zivb U994 ( .A(CUR_PERADDR_4), .Y(n1699) );
    zdffqrb CUR_PERADDR_reg_3 ( .CK(PCICLK), .D(CUR_PERADDR1050_3), .R(TRST_), 
        .Q(CUR_PERADDR_3) );
    zivb U995 ( .A(CUR_PERADDR_3), .Y(n1709) );
    zdffqrb CUR_PERADDR_reg_2 ( .CK(PCICLK), .D(CUR_PERADDR1050_2), .R(TRST_), 
        .Q(CUR_PERADDR_2) );
    zivb U996 ( .A(CUR_PERADDR_2), .Y(n1711) );
    zdffqrb CUR_PERADDR_reg_1 ( .CK(PCICLK), .D(CUR_PERADDR1050_1), .R(TRST_), 
        .Q(CUR_PERADDR_1) );
    zivb U997 ( .A(CUR_PERADDR_1), .Y(n1701) );
    zdffqrb CUR_ASYNCADDR_reg_6 ( .CK(PCICLK), .D(CUR_ASYNCADDR1138_6), .R(
        TRST_), .Q(CUR_ASYNCADDR_6) );
    zivb U998 ( .A(CUR_ASYNCADDR_6), .Y(n1706) );
    zdffqrb CUR_ASYNCADDR_reg_5 ( .CK(PCICLK), .D(CUR_ASYNCADDR1138_5), .R(
        TRST_), .Q(CUR_ASYNCADDR_5) );
    zivb U999 ( .A(CUR_ASYNCADDR_5), .Y(n1708) );
    zdffqrb CUR_ASYNCADDR_reg_4 ( .CK(PCICLK), .D(CUR_ASYNCADDR1138_4), .R(
        TRST_), .Q(CUR_ASYNCADDR_4) );
    zivb U1000 ( .A(CUR_ASYNCADDR_4), .Y(n1700) );
    zdffqrb CUR_ASYNCADDR_reg_3 ( .CK(PCICLK), .D(CUR_ASYNCADDR1138_3), .R(
        TRST_), .Q(CUR_ASYNCADDR_3) );
    zivb U1001 ( .A(CUR_ASYNCADDR_3), .Y(n1710) );
    zdffqrb CUR_ASYNCADDR_reg_2 ( .CK(PCICLK), .D(CUR_ASYNCADDR1138_2), .R(
        TRST_), .Q(CUR_ASYNCADDR_2) );
    zivb U1002 ( .A(CUR_ASYNCADDR_2), .Y(n1712) );
    zdffqrb CUR_ASYNCADDR_reg_1 ( .CK(PCICLK), .D(CUR_ASYNCADDR1138_1), .R(
        TRST_), .Q(CUR_ASYNCADDR_1) );
    zivb U1003 ( .A(CUR_ASYNCADDR_1), .Y(n1702) );
    zdffqrb SLBUI_GO_reg ( .CK(PCICLK), .D(SLBUI_GO269), .R(TRST_), .Q(
        SLBUI_GO) );
    zivb U1004 ( .A(SLBUI_GO), .Y(n1850) );
    zdffrb PERIODCMDEXE_reg ( .CK(PCICLK), .D(PERIODCMDEXE856), .R(TRST_), .Q(
        PERIODCMDEXE), .QN(SL_ERROFFSET[7]) );
    zdffqrb SLCMDSTART_reg ( .CK(PCICLK), .D(n1649), .R(TRST_), .Q(SLCMDSTART)
         );
    zdffqrb SL_PCIERR_reg ( .CK(PCICLK), .D(SL_PCIERR967), .R(TRST_), .Q(
        SL_PCIERR) );
    zdffqrb SLHCIREQ_reg ( .CK(PCICLK), .D(SLHCIREQ306), .R(TRST_), .Q(
        SLHCIREQ) );
    zdffqrb SLAVE_GO_reg ( .CK(PCICLK), .D(SLAVE_GO156), .R(TRST_), .Q(
        SLAVE_GO) );
    zivb U1005 ( .A(SLAVE_GO), .Y(n1664) );
    zdffqrb SLREAD_reg ( .CK(PCICLK), .D(SLREAD782), .R(TRST_), .Q(SLREAD) );
    zdffqrb SLAVE_ACT_reg ( .CK(PCICLK), .D(SLAVE_ACT232), .R(TRST_), .Q(
        SLAVE_ACT) );
    zdffqrb SLAVE_GO_T_reg ( .CK(PCICLK), .D(n1860), .R(TRST_), .Q(SLAVE_GO_T)
         );
    zdffqrb SLAVE_ERR_reg ( .CK(PCICLK), .D(SLAVE_ERR930), .R(TRST_), .Q(
        SLAVE_ERR) );
    zivb U1006 ( .A(SLAVE_ERR), .Y(n1688) );
    zoa21b U1007 ( .A(n1685), .B(n1724), .C(n1727), .Y(n1641) );
    znr2b U1008 ( .A(n1720), .B(n1719), .Y(n1642) );
    zaoi21b U1009 ( .A(n1661), .B(SL_ERROFFSET[7]), .C(n1747), .Y(n1643) );
    znr3d U1010 ( .A(SLBUI_GO), .B(n1742), .C(n1741), .Y(n1644) );
    zaoi21b U1011 ( .A(n1743), .B(n1744), .C(SLBUI_GO), .Y(n1645) );
    znr2b U1012 ( .A(SLBUI_GO), .B(n1676), .Y(n1646) );
    znr3d U1013 ( .A(SLBUI_GO), .B(n1745), .C(n1741), .Y(n1647) );
    zaoi21b U1014 ( .A(n1746), .B(n1744), .C(SLBUI_GO), .Y(n1648) );
    znr2b U1015 ( .A(n1851), .B(n1687), .Y(n1649) );
    zdffqrb CUR_ASYNCADDR_reg_0 ( .CK(PCICLK), .D(CUR_ASYNCADDR1138_0), .R(
        TRST_), .Q(CUR_ASYNCADDR_0) );
    zivb U1016 ( .A(CUR_ASYNCADDR_0), .Y(n1714) );
    zdffqrb CUR_PERADDR_reg_0 ( .CK(PCICLK), .D(CUR_PERADDR1050_0), .R(TRST_), 
        .Q(CUR_PERADDR_0) );
    zivb U1017 ( .A(CUR_PERADDR_0), .Y(n1713) );
    zdffqrb ASYNCADDR_reg_0 ( .CK(PCICLK), .D(ASYNCADDR465_0), .R(TRST_), .Q(
        ASYNCADDR_0) );
    zivb U1018 ( .A(ASYNCADDR_0), .Y(n1737) );
    zdffqrb PERADDR_reg_0 ( .CK(PCICLK), .D(PERADDR380_0), .R(TRST_), .Q(
        PERADDR_0) );
    zivb U1019 ( .A(PERADDR_0), .Y(n1736) );
    zivb U1020 ( .A(n1676), .Y(n1650) );
    zmux21lb U1021 ( .A(n1817), .B(n1755), .S(n1650), .Y(ASYNC_CMD_PIPE706_7)
         );
    zmux21lb U1022 ( .A(n1837), .B(n1795), .S(n1650), .Y(ASYNC_CMD_PIPE706_17)
         );
    zmux21lb U1023 ( .A(n1821), .B(n1763), .S(n1855), .Y(ASYNC_CMD_PIPE706_31)
         );
    zmux21lb U1024 ( .A(n1823), .B(n1767), .S(n1650), .Y(ASYNC_CMD_PIPE706_3)
         );
    zmux21lb U1025 ( .A(n1829), .B(n1779), .S(n1855), .Y(ASYNC_CMD_PIPE706_24)
         );
    zmux21lb U1026 ( .A(n1827), .B(n1775), .S(n1855), .Y(ASYNC_CMD_PIPE706_26)
         );
    zmux21lb U1027 ( .A(n1831), .B(n1783), .S(n1855), .Y(ASYNC_CMD_PIPE706_22)
         );
    zmux21lb U1028 ( .A(n1815), .B(n1751), .S(n1855), .Y(ASYNC_CMD_PIPE706_9)
         );
    zmux21lb U1029 ( .A(n1833), .B(n1787), .S(n1650), .Y(ASYNC_CMD_PIPE706_20)
         );
    zmux21lb U1030 ( .A(n1835), .B(n1791), .S(n1650), .Y(ASYNC_CMD_PIPE706_19)
         );
    zmux21lb U1031 ( .A(n1845), .B(n1811), .S(n1650), .Y(ASYNC_CMD_PIPE706_1)
         );
    zmux21lb U1032 ( .A(n1825), .B(n1771), .S(n1855), .Y(ASYNC_CMD_PIPE706_28)
         );
    zmux21lb U1033 ( .A(n1843), .B(n1807), .S(n1650), .Y(ASYNC_CMD_PIPE706_11)
         );
    zmux21lb U1034 ( .A(n1819), .B(n1759), .S(n1650), .Y(ASYNC_CMD_PIPE706_5)
         );
    zmux21lb U1035 ( .A(n1841), .B(n1803), .S(n1855), .Y(ASYNC_CMD_PIPE706_13)
         );
    zmux21lb U1036 ( .A(n1839), .B(n1799), .S(n1855), .Y(ASYNC_CMD_PIPE706_15)
         );
    zor2b U1037 ( .A(SLBUI_GO), .B(n1748), .Y(n1747) );
    zivb U1038 ( .A(n1676), .Y(n1748) );
    zivb U1039 ( .A(n1740), .Y(n1651) );
    zmux21lb U1040 ( .A(n1804), .B(n1805), .S(n1739), .Y(PERIOD_CMD_PIPE592_12
        ) );
    zmux21lb U1041 ( .A(n1768), .B(n1769), .S(n1739), .Y(PERIOD_CMD_PIPE592_29
        ) );
    zmux21lb U1042 ( .A(n1796), .B(n1797), .S(n1739), .Y(PERIOD_CMD_PIPE592_16
        ) );
    zmux21lb U1043 ( .A(n1800), .B(n1801), .S(n1651), .Y(PERIOD_CMD_PIPE592_14
        ) );
    zmux21lb U1044 ( .A(n1780), .B(n1781), .S(n1651), .Y(PERIOD_CMD_PIPE592_23
        ) );
    zmux21lb U1045 ( .A(n1788), .B(n1789), .S(n1651), .Y(PERIOD_CMD_PIPE592_2)
         );
    zmux21lb U1046 ( .A(n1776), .B(n1777), .S(n1651), .Y(PERIOD_CMD_PIPE592_25
        ) );
    zmux21lb U1047 ( .A(n1812), .B(n1813), .S(n1739), .Y(PERIOD_CMD_PIPE592_0)
         );
    zmux21lb U1048 ( .A(n1772), .B(n1773), .S(n1739), .Y(PERIOD_CMD_PIPE592_27
        ) );
    zmux21lb U1049 ( .A(n1784), .B(n1785), .S(n1739), .Y(PERIOD_CMD_PIPE592_21
        ) );
    zmux21lb U1050 ( .A(n1752), .B(n1753), .S(n1739), .Y(PERIOD_CMD_PIPE592_8)
         );
    zmux21lb U1051 ( .A(n1792), .B(n1793), .S(n1651), .Y(PERIOD_CMD_PIPE592_18
        ) );
    zmux21lb U1052 ( .A(n1756), .B(n1757), .S(n1651), .Y(PERIOD_CMD_PIPE592_6)
         );
    zmux21lb U1053 ( .A(n1808), .B(n1809), .S(n1739), .Y(PERIOD_CMD_PIPE592_10
        ) );
    zmux21lb U1054 ( .A(n1760), .B(n1761), .S(n1651), .Y(PERIOD_CMD_PIPE592_4)
         );
    zmux21lb U1055 ( .A(n1764), .B(n1765), .S(n1651), .Y(PERIOD_CMD_PIPE592_30
        ) );
    zao22b U1056 ( .A(n1857), .B(PERIOD_PIPE_1), .C(n1661), .D(PERIODCMDEXE), 
        .Y(n1852) );
    zor2b U1057 ( .A(SLADDR[7]), .B(n1719), .Y(n1740) );
    zivb U1058 ( .A(n1740), .Y(n1857) );
    zor3b U1059 ( .A(SLSM_2), .B(SLSM_0), .C(n1652), .Y(SLADDR[7]) );
    zao211b U1060 ( .A(SLSM_1), .B(n1654), .C(n1655), .D(n1656), .Y(
        SLHCIREQ306) );
    zoa21d U1061 ( .A(SLAVE_ACT), .B(EHCI_MAC_EOT), .C(SLAVEMODE), .Y(
        SLAVE_GO156) );
    zan4b U1062 ( .A(n1657), .B(n1652), .C(n1654), .D(n1641), .Y(SLBUI_GO269)
         );
    zoa21d U1063 ( .A(n1658), .B(n1649), .C(SLAVEMODE), .Y(SLAVE_ACT232) );
    zao222b U1064 ( .A(n1646), .B(n1659), .C(n1660), .D(n1661), .E(n1643), .F(
        ASYNC_PIPE_0), .Y(ASYNC_PIPE668_0) );
    zao222b U1065 ( .A(n1666), .B(n1667), .C(n1668), .D(n1661), .E(
        PERIOD_PIPE_0), .F(n1669), .Y(PERIOD_PIPE554_0) );
    zoa21d U1066 ( .A(n1675), .B(n1676), .C(n1677), .Y(n1674) );
    zoa21d U1067 ( .A(PERIODCMDEXE), .B(n1657), .C(EHCI_MAC_EOT), .Y(n1682) );
    zoa21d U1068 ( .A(n1683), .B(n1686), .C(n1652), .Y(n1685) );
    zoa21d U1069 ( .A(n1641), .B(SLSMNXT_1), .C(n1687), .Y(n1656) );
    zan4b U1070 ( .A(CUR_PERADDR_2), .B(CUR_PERADDR_3), .C(CUR_PERADDR_0), .D(
        n1690), .Y(n1689) );
    zan4b U1071 ( .A(CUR_ASYNCADDR_2), .B(CUR_ASYNCADDR_3), .C(CUR_ASYNCADDR_0
        ), .D(n1692), .Y(n1691) );
    zor3b U1072 ( .A(n1652), .B(n1722), .C(n1719), .Y(n1676) );
    zor3b U1073 ( .A(GEN_PERR), .B(SLAVE_ERR), .C(n1704), .Y(n1694) );
    zor6b U1074 ( .A(PIDERR), .B(SL_DATA_PIDERR), .C(CRCERR), .D(SL_ACK_ERR), 
        .E(SL_ET_ERR), .F(SL_SE_ERR), .Y(n1848) );
    zcx8d U1075 ( .A(n1849), .B(n1716), .C(ASYNC_FULL), .D(n1725), .E(n1642), 
        .Y(n1677) );
    zcx8d U1076 ( .A(SLADDR[7]), .B(n1642), .C(n1655), .D(n1652), .E(TDMAEND), 
        .Y(n1679) );
    zan4b U1077 ( .A(CUR_PERADDR_5), .B(CUR_PERADDR_6), .C(CUR_PERADDR_1), .D(
        CUR_PERADDR_4), .Y(n1690) );
    zan4b U1078 ( .A(CUR_ASYNCADDR_5), .B(CUR_ASYNCADDR_6), .C(CUR_ASYNCADDR_1
        ), .D(CUR_ASYNCADDR_4), .Y(n1692) );
    zbfb U1079 ( .A(SLAVE_GO), .Y(n1860) );
endmodule


module TESTPKTCTL ( PCICLK, TRST_, TEST_PACKET, RUN, EHCI_MAC_EOT, TESTPKTOK, 
    TBUI_GO, TCMDSTART );
input  PCICLK, TRST_, TEST_PACKET, RUN, EHCI_MAC_EOT, TESTPKTOK;
output TBUI_GO, TCMDSTART;
    wire TEST_START, SPAREO6, SPAREO0_, TCMDST, SPAREO8, SPAREO1, SPAREO9, 
        SPAREO0, TCMDST_T, SPAREO7, SPAREO5, TEST_START_T, SPAREO2, SPAREO1_, 
        SPAREO3, TEST_START69, SPAREO4, n155, n156, n157, n158, n159;
    zdffrb SPARE600 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE607 ( .A(SPAREO4), .Y(SPAREO5) );
    znd3b SPARE609 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE601 ( .CK(1'b0), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE608 ( .A(SPAREO5), .Y(SPAREO6) );
    znr3b SPARE606 ( .A(SPAREO2), .B(TEST_START_T), .C(SPAREO0_), .Y(SPAREO4)
         );
    zaoi211b SPARE603 ( .A(SPAREO4), .B(TEST_START), .C(SPAREO6), .D(1'b0), 
        .Y(SPAREO8) );
    zoai21b SPARE604 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE602 ( .A(SPAREO0), .B(TCMDST), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE605 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zan2b U41 ( .A(n155), .B(TEST_PACKET), .Y(TEST_START69) );
    zdffqrb TCMDST_reg ( .CK(PCICLK), .D(TESTPKTOK), .R(TRST_), .Q(TCMDST) );
    zdffqrb TEST_START_T_reg ( .CK(PCICLK), .D(n159), .R(TRST_), .Q(
        TEST_START_T) );
    zdffqrb TEST_START_reg ( .CK(PCICLK), .D(TEST_START69), .R(TRST_), .Q(
        TEST_START) );
    zdffqrb TCMDST_T_reg ( .CK(PCICLK), .D(n157), .R(TRST_), .Q(TCMDST_T) );
    zinr2b U42 ( .A(TESTPKTOK), .B(TCMDST_T), .Y(TCMDSTART) );
    zinr2b U43 ( .A(TEST_START), .B(TEST_START_T), .Y(TBUI_GO) );
    zinr2b U44 ( .A(EHCI_MAC_EOT), .B(RUN), .Y(n155) );
    zivb U45 ( .A(TCMDST), .Y(n156) );
    zivb U46 ( .A(n156), .Y(n157) );
    zivb U47 ( .A(TEST_START), .Y(n158) );
    zivb U48 ( .A(n158), .Y(n159) );
endmodule


module DBGCTL ( EN_DBG_PORT, GEN_PERR, DBGPORT_SC, DBGPORT_PID, DBGPORT_ADDR, 
    DBG_COMPL, DBG_XACTERR, DBG_RXPID, DBG_RXBCNT, DBG_CMDSTART_REQ, TRAN_CMD, 
    DBG_ACT, DBG_CMDSTART, EHCI_MAC_EOT, CRCERR, BABBLE, PIDERR, TMOUT, RXACK, 
    RXPID, RXBCNT, PCICLK, TRST_ );
input  [31:0] DBGPORT_SC;
output [7:0] DBG_RXPID;
output [3:0] DBG_RXBCNT;
input  [7:0] RXPID;
input  [31:0] DBGPORT_PID;
input  [31:0] DBGPORT_ADDR;
output [51:0] TRAN_CMD;
input  [10:0] RXBCNT;
input  EN_DBG_PORT, GEN_PERR, DBG_CMDSTART, EHCI_MAC_EOT, CRCERR, BABBLE, 
    PIDERR, TMOUT, RXACK, PCICLK, TRST_;
output DBG_COMPL, DBG_XACTERR, DBG_CMDSTART_REQ, DBG_ACT;
    wire DBG_RXBCNT303_3, DBGSMNXT_3, SPAREO6, DBGSM_2, SPAREO0_, RX_PID265_2, 
        DBG_CMDSTART_P, SPAREO1, DBG_CMDSTART_EOT341, RX_PID265_3, SPAREO9, 
        DBG_GO_T, SPAREO0, DBGSMNXT_2, SPAREO7, DBG_RXBCNT303_2, DBGSM_3, 
        DBG_XACTERR228, DBG_RXBCNT303_0, SPAREO5, DBGSMNXT_0, DBGSM_1, 
        RX_PID265_1, SPAREO2, DBG_GO_2T, RX_PID265_0, SPAREO3, SPAREO1_, 
        DBG_CMDSTART_EOT, n550, SPAREO4, DBGSMNXT_1, DBG_RXBCNT303_1, DBGSM_0, 
        n501, n502, n503, n504, n525, n526, n527, n528, n529, n530, n531, n532, 
        n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
        n545, n546, n547, n548, n551, n552, n553;
    assign TRAN_CMD[51] = 1'b0;
    assign TRAN_CMD[50] = 1'b0;
    assign TRAN_CMD[49] = 1'b0;
    assign TRAN_CMD[48] = 1'b0;
    assign TRAN_CMD[47] = 1'b0;
    assign TRAN_CMD[46] = 1'b0;
    assign TRAN_CMD[45] = 1'b0;
    assign TRAN_CMD[44] = 1'b0;
    assign TRAN_CMD[28] = 1'b0;
    assign TRAN_CMD[27] = 1'b0;
    assign TRAN_CMD[26] = 1'b0;
    assign TRAN_CMD[25] = 1'b0;
    assign TRAN_CMD[24] = 1'b0;
    assign TRAN_CMD[23] = 1'b0;
    assign TRAN_CMD[22] = 1'b0;
    assign TRAN_CMD[21] = 1'b0;
    assign TRAN_CMD[20] = 1'b0;
    assign TRAN_CMD[19] = 1'b0;
    assign TRAN_CMD[18] = 1'b0;
    assign TRAN_CMD[17] = 1'b0;
    assign TRAN_CMD[16] = 1'b0;
    assign TRAN_CMD[15] = 1'b0;
    assign TRAN_CMD[14] = 1'b0;
    assign TRAN_CMD[13] = 1'b0;
    assign TRAN_CMD[12] = 1'b0;
    assign TRAN_CMD[11] = 1'b0;
    assign TRAN_CMD[10] = 1'b0;
    assign TRAN_CMD[7] = 1'b0;
    assign TRAN_CMD[6] = 1'b0;
    assign TRAN_CMD[5] = 1'b0;
    assign TRAN_CMD[4] = 1'b1;
    assign TRAN_CMD[0] = 1'b0;
    zoai21b SPARE_DBGC5 ( .A(SPAREO1), .B(DBG_GO_T), .C(SPAREO9), .Y(SPAREO3)
         );
    zaoi211b SPARE_DBGC2 ( .A(SPAREO0), .B(DBG_GO_2T), .C(SPAREO1_), .D(1'b0), 
        .Y(SPAREO2) );
    zaoi211b SPARE_DBGC3 ( .A(SPAREO4), .B(DBG_CMDSTART_P), .C(SPAREO6), .D(
        1'b0) );
    zoai21b SPARE_DBGC4 ( .A(SPAREO0), .B(n550), .C(1'b0), .Y(SPAREO9) );
    znr3b SPARE_DBGC6 ( .A(SPAREO2), .B(n501), .C(SPAREO0_), .Y(SPAREO4) );
    zdffrb SPARE_DBGC1 ( .CK(PCICLK), .D(SPAREO7), .R(TRST_), .Q(SPAREO1), 
        .QN(SPAREO1_) );
    zivb SPARE_DBGC8 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE_DBGC0 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE_DBGC9 ( .A(SPAREO3), .B(SPAREO6), .C(1'b0), .Y(SPAREO7) );
    zivb SPARE_DBGC7 ( .A(SPAREO4), .Y(SPAREO5) );
    zan2b U146 ( .A(n504), .B(n538), .Y(n537) );
    zan2b U147 ( .A(DBGSM_2), .B(DBGSM_3), .Y(n539) );
    zor2b U148 ( .A(DBGSM_2), .B(n540), .Y(n541) );
    zor2b U149 ( .A(DBGSM_3), .B(DBGSM_2), .Y(n545) );
    zmux21hb U150 ( .A(DBG_RXPID[3]), .B(RXPID[3]), .S(n501), .Y(RX_PID265_3)
         );
    zmux21hb U151 ( .A(DBG_RXPID[2]), .B(RXPID[2]), .S(n501), .Y(RX_PID265_2)
         );
    zmux21hb U152 ( .A(DBG_RXPID[1]), .B(RXPID[1]), .S(n501), .Y(RX_PID265_1)
         );
    zmux21hb U153 ( .A(DBG_RXPID[0]), .B(RXPID[0]), .S(n501), .Y(RX_PID265_0)
         );
    zmux21hb U154 ( .A(DBG_RXBCNT[3]), .B(RXBCNT[3]), .S(n501), .Y(
        DBG_RXBCNT303_3) );
    zmux21hb U155 ( .A(DBG_RXBCNT[2]), .B(RXBCNT[2]), .S(n501), .Y(
        DBG_RXBCNT303_2) );
    zmux21hb U156 ( .A(DBG_RXBCNT[1]), .B(RXBCNT[1]), .S(n501), .Y(
        DBG_RXBCNT303_1) );
    zmux21hb U157 ( .A(DBG_RXBCNT[0]), .B(RXBCNT[0]), .S(n501), .Y(
        DBG_RXBCNT303_0) );
    zmux21lb U158 ( .A(n527), .B(n537), .S(DBGSM_0), .Y(n531) );
    zao21b U159 ( .A(n503), .B(n529), .C(n532), .Y(DBGSMNXT_1) );
    zivb U160 ( .A(GEN_PERR), .Y(n535) );
    zao22b U161 ( .A(DBG_CMDSTART), .B(n502), .C(n525), .D(n526), .Y(
        DBGSMNXT_3) );
    zivb U162 ( .A(n543), .Y(n525) );
    zor2b U163 ( .A(DBG_CMDSTART), .B(n529), .Y(n526) );
    zivb U164 ( .A(EHCI_MAC_EOT), .Y(n529) );
    zao22b U165 ( .A(n502), .B(n533), .C(n503), .D(EHCI_MAC_EOT), .Y(
        DBGSMNXT_2) );
    zivb U166 ( .A(DBG_CMDSTART), .Y(n533) );
    zmux21hb U167 ( .A(DBG_XACTERR), .B(n548), .S(n501), .Y(DBG_XACTERR228) );
    zor2b U168 ( .A(DBG_COMPL), .B(n527), .Y(DBG_ACT) );
    zor2b U169 ( .A(DBGSM_1), .B(n545), .Y(n527) );
    zivb U170 ( .A(DBG_ACT), .Y(n536) );
    zivb U171 ( .A(n527), .Y(n538) );
    zivb U172 ( .A(DBGPORT_SC[4]), .Y(TRAN_CMD[1]) );
    zivb U173 ( .A(DBGPORT_SC[4]), .Y(TRAN_CMD[3]) );
    zan2b U174 ( .A(DBG_CMDSTART_P), .B(n528), .Y(DBG_CMDSTART_REQ) );
    zor2b U175 ( .A(DBGSMNXT_3), .B(DBGSM_2), .Y(DBG_CMDSTART_P) );
    zdffrb RX_PID_reg_3 ( .CK(PCICLK), .D(RX_PID265_3), .R(TRST_), .Q(
        DBG_RXPID[3]), .QN(DBG_RXPID[7]) );
    zdffrb RX_PID_reg_2 ( .CK(PCICLK), .D(RX_PID265_2), .R(TRST_), .Q(
        DBG_RXPID[2]), .QN(DBG_RXPID[6]) );
    zdffrb RX_PID_reg_1 ( .CK(PCICLK), .D(RX_PID265_1), .R(TRST_), .Q(
        DBG_RXPID[1]), .QN(DBG_RXPID[5]) );
    zdffrb RX_PID_reg_0 ( .CK(PCICLK), .D(RX_PID265_0), .R(TRST_), .Q(
        DBG_RXPID[0]), .QN(DBG_RXPID[4]) );
    zdffqrb DBG_RXBCNT_reg_3 ( .CK(PCICLK), .D(DBG_RXBCNT303_3), .R(TRST_), 
        .Q(DBG_RXBCNT[3]) );
    zdffqrb DBG_RXBCNT_reg_2 ( .CK(PCICLK), .D(DBG_RXBCNT303_2), .R(TRST_), 
        .Q(DBG_RXBCNT[2]) );
    zdffqrb DBG_RXBCNT_reg_1 ( .CK(PCICLK), .D(DBG_RXBCNT303_1), .R(TRST_), 
        .Q(DBG_RXBCNT[1]) );
    zdffqrb DBG_RXBCNT_reg_0 ( .CK(PCICLK), .D(DBG_RXBCNT303_0), .R(TRST_), 
        .Q(DBG_RXBCNT[0]) );
    zdffqrb DBG_CMDSTART_EOT_reg ( .CK(PCICLK), .D(n553), .R(TRST_), .Q(
        DBG_CMDSTART_EOT) );
    zivb U176 ( .A(DBG_CMDSTART_EOT), .Y(n528) );
    zdffqrb DBG_GO_2T_reg ( .CK(PCICLK), .D(n552), .R(TRST_), .Q(DBG_GO_2T) );
    zdffqrb DBG_GO_T_reg ( .CK(PCICLK), .D(DBGPORT_SC[5]), .R(TRST_), .Q(
        DBG_GO_T) );
    zdffqsb DBGSM_reg_0 ( .CK(PCICLK), .D(DBGSMNXT_0), .S(TRST_), .Q(DBGSM_0)
         );
    zdffqrb DBGSM_reg_1 ( .CK(PCICLK), .D(DBGSMNXT_1), .R(TRST_), .Q(DBGSM_1)
         );
    zivb U177 ( .A(DBGSM_1), .Y(n546) );
    zdffqrb DBGSM_reg_4 ( .CK(PCICLK), .D(n501), .R(TRST_), .Q(DBG_COMPL) );
    zdffqrb DBGSM_reg_3 ( .CK(PCICLK), .D(DBGSMNXT_3), .R(TRST_), .Q(DBGSM_3)
         );
    zivb U178 ( .A(DBGSM_3), .Y(n542) );
    zdffqrb DBGSM_reg_2 ( .CK(PCICLK), .D(DBGSMNXT_2), .R(TRST_), .Q(DBGSM_2)
         );
    zivb U179 ( .A(DBGSM_2), .Y(n544) );
    zdffqrb DBG_XACTERR_reg ( .CK(PCICLK), .D(DBG_XACTERR228), .R(TRST_), .Q(
        DBG_XACTERR) );
    znr2d U180 ( .A(n526), .B(n543), .Y(n501) );
    znr4b U181 ( .A(DBGSM_3), .B(DBGSM_1), .C(n544), .D(n540), .Y(n502) );
    znr3b U182 ( .A(DBGSM_3), .B(n546), .C(n541), .Y(n503) );
    zan2b U183 ( .A(n547), .B(EN_DBG_PORT), .Y(n504) );
    zivb U184 ( .A(DBGPORT_SC[4]), .Y(n550) );
    ziv11b U185 ( .A(DBGPORT_SC[4]), .Y(TRAN_CMD[2]), .Z(TRAN_CMD[8]) );
    zivb U186 ( .A(DBGPORT_SC[4]), .Y(TRAN_CMD[9]) );
    zbfb U187 ( .A(DBGPORT_ADDR[0]), .Y(TRAN_CMD[29]) );
    zbfb U188 ( .A(DBGPORT_ADDR[1]), .Y(TRAN_CMD[30]) );
    zbfb U189 ( .A(DBGPORT_ADDR[2]), .Y(TRAN_CMD[31]) );
    zbfb U190 ( .A(DBGPORT_ADDR[3]), .Y(TRAN_CMD[32]) );
    zbfb U191 ( .A(DBGPORT_ADDR[8]), .Y(TRAN_CMD[33]) );
    zbfb U192 ( .A(DBGPORT_ADDR[9]), .Y(TRAN_CMD[34]) );
    zbfb U193 ( .A(DBGPORT_ADDR[10]), .Y(TRAN_CMD[35]) );
    zbfb U194 ( .A(DBGPORT_ADDR[11]), .Y(TRAN_CMD[36]) );
    zbfb U195 ( .A(DBGPORT_ADDR[12]), .Y(TRAN_CMD[37]) );
    zbfb U196 ( .A(DBGPORT_ADDR[13]), .Y(TRAN_CMD[38]) );
    zbfb U197 ( .A(DBGPORT_ADDR[14]), .Y(TRAN_CMD[39]) );
    zbfb U198 ( .A(DBGPORT_SC[0]), .Y(TRAN_CMD[40]) );
    zbfb U199 ( .A(DBGPORT_SC[1]), .Y(TRAN_CMD[41]) );
    zbfb U200 ( .A(DBGPORT_SC[2]), .Y(TRAN_CMD[42]) );
    zbfb U201 ( .A(DBGPORT_SC[3]), .Y(TRAN_CMD[43]) );
    zoa21d U202 ( .A(DBG_CMDSTART), .B(DBG_CMDSTART_EOT), .C(n529), .Y(
        DBG_CMDSTART_EOT341) );
    zor3b U203 ( .A(GEN_PERR), .B(n530), .C(n531), .Y(DBGSMNXT_0) );
    zinr2b U204 ( .A(DBGPORT_SC[4]), .B(RXACK), .Y(n534) );
    zan4b U205 ( .A(DBGSM_0), .B(n504), .C(n535), .D(n536), .Y(n532) );
    zor3b U206 ( .A(DBG_COMPL), .B(DBGSM_0), .C(GEN_PERR), .Y(n540) );
    zor3b U207 ( .A(DBGSM_1), .B(n542), .C(n541), .Y(n543) );
    zor5b U208 ( .A(TMOUT), .B(PIDERR), .C(BABBLE), .D(CRCERR), .E(n534), .Y(
        n548) );
    zinr2b U209 ( .A(DBG_GO_T), .B(DBG_GO_2T), .Y(n547) );
    zao211b U210 ( .A(DBGSM_1), .B(n545), .C(DBG_COMPL), .D(n539), .Y(n530) );
    zivb U211 ( .A(DBG_GO_T), .Y(n551) );
    zivb U212 ( .A(n551), .Y(n552) );
    zbfb U213 ( .A(DBG_CMDSTART_EOT341), .Y(n553) );
endmodule


module DBG_FMTIMER ( EN_DBG_PORT, DBG_OWNER, DBG_ENABLE, RUN, EHCI_SOFGEN, 
    DBG_SOFGEN, SOFGEN, EHCI_DBG_RUN, MAC_EOT, EHCI_DBG_MAC_EOT, PRESOF, 
    EHCI_DBG_PRESOF, EHCI_EOF1, EOF1, CLK60M, TRST_ );
input  EN_DBG_PORT, DBG_OWNER, DBG_ENABLE, RUN, EHCI_SOFGEN, MAC_EOT, PRESOF, 
    EHCI_EOF1, CLK60M, TRST_;
output DBG_SOFGEN, SOFGEN, EHCI_DBG_RUN, EHCI_DBG_MAC_EOT, EHCI_DBG_PRESOF, 
    EOF1;
    wire SPAREO6, DBG_FMREMN131_2, DBG_FMREMN_4, DBG_FMREMN121_3, 
        DBG_FMREMN121_4, DBG_FMREMN_3, SPAREO0_, SPAREO8, DBG_FMREMN131_5, 
        DBG_MACEOT_MASK209, SPAREO1, SPAREO9, DBG_FMREMN131_4, DBG_FMREMN121_5, 
        DBG_FMREMN_2, SPAREO0, SPAREO7, DBG_FMREMN_5, DBG_FMREMN121_2, 
        DBG_TIMER_EN, DBG_FMREMN131_3, DBG_SOFGEN172, SPAREO5, DBG_FMREMN131_8, 
        DBG_FMREMN131_1, DBG_FMREMN_7, DBG_FMREMN_0, DBG_FMREMN121_0, 
        DBG_FMREMN121_7, DBG_MACEOT_MASK, DBG_FMREMN131_6, RUN_CLK60M, SPAREO2, 
        DBG_AND, DBG_FMREMN131_7, DBG_FMREMN_1, DBG_FMREMN121_6, SPAREO3, 
        SPAREO1_, DBG_FMREMN_8, DBG_FMREMN121_8, SPAREO4, DBG_FMREMN_6, 
        DBG_FMREMN121_1, DBG_FMREMN131_0, add_32_carry_8, add_32_carry_6, 
        add_32_carry_7, add_32_carry_2, add_32_carry_5, add_32_carry_4, 
        add_32_carry_3, n394, n395, n396, n397, n398;
    zoai21b SPARE_DBGTM5 ( .A(SPAREO1), .B(RUN_CLK60M), .C(SPAREO9), .Y(
        SPAREO3) );
    zaoi211b SPARE_DBGTM2 ( .A(SPAREO0), .B(DBG_SOFGEN), .C(SPAREO1_), .D(1'b0
        ), .Y(SPAREO2) );
    zaoi211b SPARE_DBGTM3 ( .A(SPAREO4), .B(DBG_TIMER_EN), .C(SPAREO6), .D(
        1'b0), .Y(SPAREO8) );
    zoai21b SPARE_DBGTM4 ( .A(SPAREO0), .B(SPAREO8), .C(DBG_MACEOT_MASK), .Y(
        SPAREO9) );
    znr3b SPARE_DBGTM6 ( .A(SPAREO2), .B(DBG_AND), .C(SPAREO0_), .Y(SPAREO4)
         );
    zdffrb SPARE_DBGTM1 ( .CK(CLK60M), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), 
        .QN(SPAREO1_) );
    zdffrb SPARE_DBGTM0 ( .CK(CLK60M), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE_DBGTM8 ( .A(SPAREO5), .Y(SPAREO6) );
    znd3b SPARE_DBGTM9 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb SPARE_DBGTM7 ( .A(SPAREO4), .Y(SPAREO5) );
    zan2b U101 ( .A(DBG_FMREMN121_8), .B(DBG_TIMER_EN), .Y(DBG_FMREMN131_8) );
    zan2b U102 ( .A(DBG_FMREMN121_7), .B(DBG_TIMER_EN), .Y(DBG_FMREMN131_7) );
    zhadrb add_32_U1_1_7 ( .A(DBG_FMREMN_7), .B(add_32_carry_7), .CO(
        add_32_carry_8), .S(DBG_FMREMN121_7) );
    zan2b U103 ( .A(DBG_FMREMN121_6), .B(DBG_TIMER_EN), .Y(DBG_FMREMN131_6) );
    zhadrb add_32_U1_1_6 ( .A(DBG_FMREMN_6), .B(add_32_carry_6), .CO(
        add_32_carry_7), .S(DBG_FMREMN121_6) );
    zan2b U104 ( .A(DBG_FMREMN121_5), .B(DBG_TIMER_EN), .Y(DBG_FMREMN131_5) );
    zhadrb add_32_U1_1_5 ( .A(DBG_FMREMN_5), .B(add_32_carry_5), .CO(
        add_32_carry_6), .S(DBG_FMREMN121_5) );
    zan2b U105 ( .A(DBG_FMREMN121_4), .B(DBG_TIMER_EN), .Y(DBG_FMREMN131_4) );
    zhadrb add_32_U1_1_4 ( .A(DBG_FMREMN_4), .B(add_32_carry_4), .CO(
        add_32_carry_5), .S(DBG_FMREMN121_4) );
    zan2b U106 ( .A(DBG_FMREMN121_3), .B(DBG_TIMER_EN), .Y(DBG_FMREMN131_3) );
    zhadrb add_32_U1_1_3 ( .A(DBG_FMREMN_3), .B(add_32_carry_3), .CO(
        add_32_carry_4), .S(DBG_FMREMN121_3) );
    zan2b U107 ( .A(DBG_FMREMN121_2), .B(DBG_TIMER_EN), .Y(DBG_FMREMN131_2) );
    zhadrb add_32_U1_1_2 ( .A(DBG_FMREMN_2), .B(add_32_carry_2), .CO(
        add_32_carry_3), .S(DBG_FMREMN121_2) );
    zan2b U108 ( .A(DBG_FMREMN121_1), .B(DBG_TIMER_EN), .Y(DBG_FMREMN131_1) );
    zhadrb add_32_U1_1_1 ( .A(DBG_FMREMN_1), .B(DBG_FMREMN_0), .CO(
        add_32_carry_2), .S(DBG_FMREMN121_1) );
    zan2b U109 ( .A(DBG_FMREMN121_0), .B(DBG_TIMER_EN), .Y(DBG_FMREMN131_0) );
    zan2b U110 ( .A(DBG_FMREMN_3), .B(DBG_FMREMN_5), .Y(n394) );
    zivb U111 ( .A(MAC_EOT), .Y(n395) );
    zan2b U112 ( .A(EHCI_EOF1), .B(n396), .Y(EOF1) );
    zan2b U113 ( .A(PRESOF), .B(n396), .Y(EHCI_DBG_PRESOF) );
    zor2b U114 ( .A(DBG_AND), .B(RUN), .Y(EHCI_DBG_RUN) );
    zivb U115 ( .A(n398), .Y(DBG_AND) );
    znd3b U116 ( .A(DBG_OWNER), .B(DBG_ENABLE), .C(EN_DBG_PORT), .Y(n398) );
    zmux21hb U117 ( .A(EHCI_SOFGEN), .B(DBG_SOFGEN), .S(DBG_TIMER_EN), .Y(
        SOFGEN) );
    zivb U118 ( .A(n396), .Y(DBG_TIMER_EN) );
    zor2b U119 ( .A(RUN_CLK60M), .B(n398), .Y(n396) );
    zdffqrb DBG_FMREMN_reg_8 ( .CK(CLK60M), .D(DBG_FMREMN131_8), .R(TRST_), 
        .Q(DBG_FMREMN_8) );
    zdffqrb DBG_FMREMN_reg_7 ( .CK(CLK60M), .D(DBG_FMREMN131_7), .R(TRST_), 
        .Q(DBG_FMREMN_7) );
    zdffqrb DBG_FMREMN_reg_6 ( .CK(CLK60M), .D(DBG_FMREMN131_6), .R(TRST_), 
        .Q(DBG_FMREMN_6) );
    zdffqrb DBG_FMREMN_reg_5 ( .CK(CLK60M), .D(DBG_FMREMN131_5), .R(TRST_), 
        .Q(DBG_FMREMN_5) );
    zdffqrb DBG_FMREMN_reg_4 ( .CK(CLK60M), .D(DBG_FMREMN131_4), .R(TRST_), 
        .Q(DBG_FMREMN_4) );
    zdffqrb DBG_FMREMN_reg_3 ( .CK(CLK60M), .D(DBG_FMREMN131_3), .R(TRST_), 
        .Q(DBG_FMREMN_3) );
    zdffqrb DBG_FMREMN_reg_2 ( .CK(CLK60M), .D(DBG_FMREMN131_2), .R(TRST_), 
        .Q(DBG_FMREMN_2) );
    zdffqrb DBG_FMREMN_reg_1 ( .CK(CLK60M), .D(DBG_FMREMN131_1), .R(TRST_), 
        .Q(DBG_FMREMN_1) );
    zdffqrb DBG_FMREMN_reg_0 ( .CK(CLK60M), .D(DBG_FMREMN131_0), .R(TRST_), 
        .Q(DBG_FMREMN_0) );
    zivb U120 ( .A(DBG_FMREMN_0), .Y(DBG_FMREMN121_0) );
    zdffqrb DBG_SOFGEN_reg ( .CK(CLK60M), .D(DBG_SOFGEN172), .R(TRST_), .Q(
        DBG_SOFGEN) );
    zdffqb RUN_CLK60M_reg ( .CK(CLK60M), .D(RUN), .Q(RUN_CLK60M) );
    zdffqsb DBG_MACEOT_MASK_reg ( .CK(CLK60M), .D(DBG_MACEOT_MASK209), .S(
        TRST_), .Q(DBG_MACEOT_MASK) );
    zivb U121 ( .A(DBG_MACEOT_MASK), .Y(n397) );
    zxo2b U122 ( .A(add_32_carry_8), .B(DBG_FMREMN_8), .Y(DBG_FMREMN121_8) );
    zan8b U123 ( .A(DBG_FMREMN_6), .B(DBG_FMREMN_8), .C(DBG_FMREMN_7), .D(n394
        ), .E(DBG_FMREMN_1), .F(DBG_FMREMN_4), .G(DBG_FMREMN_2), .H(
        DBG_FMREMN_0), .Y(DBG_SOFGEN172) );
    zao21b U124 ( .A(DBG_MACEOT_MASK), .B(n395), .C(RUN_CLK60M), .Y(
        DBG_MACEOT_MASK209) );
    zao21b U125 ( .A(EN_DBG_PORT), .B(n397), .C(MAC_EOT), .Y(EHCI_DBG_MAC_EOT)
         );
endmodule

// USB 2.0 EHCI control module

module EHCI ( PCI1WAIT, HCIMRDY1, HCIMRDY2, RDYACK, HCICOMPL1, HCICOMPL2,
              MABORTS, TABORTR, HCIGNT1, HCIGNT2, /*PCICLK,*/ TRST_,
              PAROPT, PERRS, SERRS, PMSTR1, PMSTR3, MADDR1, MADDR3, ADI, SADI,
	      ASYNC_EN, PERIOD_EN, SOFGEN, EOFTERM, FEMPTY1, FEMPTY2,
	      FEMPTY3, FEMPTY4,
	      EHCIREQ1, EHCIREQ2, SLHCIREQ, CLK60M, FLADJ, REDUCE, EOF1, EOF2,
	      FRNUM, SOFV, WR_FRNUM, FRLSTSIZE, FRNUM_PCLK_LATCH,
	      RUN, HCHALT, FLBASE, HCIADR1, HCIADR2, CMDSTART, MAC_EOT, TXSOF,
	      BUI_GO1, BUI_GO2, BUI_GO3, BUI_GO4, TDMAEND1,
	      TDMAEND2, TDMAEND3, TDMAEND4, /*TXTHRESH,*/
	      EOT1, EOT2, EOT3, EOT4,
	      CRCERR, RXERR1, RXERR2, RXERR3, RXERR4, ACTLEN, BABBLE,
	      HCIADD1, HCIADD2, HCIMWR1, HCIMWR2, /*BOUNDRY,*/ WPR1, WPR2,
	      PIDERR, ASYNCLISTADDR, RECLAMATION, TMOUT, RXNAK, RXNYET, RXSTALL,
	      RXACK, RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXPIDERR, RXPID,
	      TOGMATCH, SPD, ASYNC_ACT, PERIOD_ACT, RUN_C, WR_ASYNCADDR,
	      TRAN_CMD1, TRAN_CMD2, TRAN_CMD3, TRAN_CMD4, MAXLEN,
	      CREQ1, CREQ2, CREQ3, CREQ4, PCIDMA_SEL, USBDMA_SEL,
	      RXBCNT, ROLLOVER_S,
	      EN_DBG_PORT, DBGPORT_SC, DBGPORT_PID, DBGPORT_ADDR,
	      DBG_COMPL, DBG_XACTERR, DBG_RXPID, DBG_RXBCNT, DBG_TRAN_CMD,
	      DBG_SEL, EHCI_DBG_MAC_EOT, DBG_IDLE,
	      INTTHRESHOLD, USBINT, USBINT_S, ERRINT, ERRINT_S, /*IOCSPDINT,
	      USBERRINT,*/ USBINT_EN, ERRINT_EN, INTDOORBELL, INTASYNC_EN,
	      INTASYNC_S, INTASYNC, ASYNCINT, EHCIEXE, TEST_PACKET,
	      TESTPKTOK, SWDBG, HSERR_S, SLAVEMODE, SLAVE_ACT,
	      BMUCRST_, SLADDR, SLREAD, DATARDY, MDO,
	      PERIOD_CMD, ASYNC_CMD, SL_PERIOD, SL_ERROFFSET,
	      SL_DATA_PIDERR, SL_ET_ERR, SL_SE_ERR, SL_ACK_ERR,
	      SL_PCIERR, SLAVE_ERR,
	      EHCI_IDLE, TD_IDLE1, TD_IDLE2, TD_IDLE3, TD_IDLE4,
	      TD_PARSE_GO1, TD_PARSE_GO2, TD_PARSE_GO3, TD_PARSE_GO4,
	      EHCIFLOW_PCLK, EHCI_DMA1_PCLK, EHCI_DMA2_PCLK,
	      EHCI_DMA3_PCLK, EHCI_DMA4_PCLK,
	      EHCIFLOW_CACHE_PCLK, EHCI_DMA1_CACHE_PCLK, EHCI_DMA2_CACHE_PCLK,
	      EHCI_DMA3_CACHE_PCLK, EHCI_DMA4_CACHE_PCLK, DBG_PCLK,
	      UGNTI1_, UGNTI3_, SLEEPTIME_SEL, ATPG_ENI
            );
input	DBG_PCLK;
output	DBG_IDLE;
output	FRNUM_PCLK_LATCH;
input	SLEEPTIME_SEL;	// option to reduce EHCI sleep time
input   EHCIFLOW_PCLK, EHCI_DMA1_PCLK, EHCI_DMA2_PCLK,
	EHCI_DMA3_PCLK, EHCI_DMA4_PCLK;
input   EHCIFLOW_CACHE_PCLK, EHCI_DMA1_CACHE_PCLK, EHCI_DMA2_CACHE_PCLK,
	EHCI_DMA3_CACHE_PCLK, EHCI_DMA4_CACHE_PCLK;
input   PCI1WAIT, RDYACK, MABORTS, TABORTR, PAROPT, PERRS, SERRS,
	PMSTR1, PMSTR3;
//input	MADDR1, MADDR3;
output	MADDR1, MADDR3;
input	UGNTI1_, UGNTI3_;
output  HCICOMPL1, HCICOMPL2, HCIMRDY1, HCIMRDY2;
input   /*PCICLK,*/ TRST_, HCIGNT1, HCIGNT2;
input	[31:0]	ADI;		// data bus to latch data
input	[31:0]	SADI;		// slave data path
input	ASYNC_EN, PERIOD_EN, EOFTERM;
output	EHCIREQ1, EHCIREQ2, SLHCIREQ;
input	CLK60M, REDUCE, WR_FRNUM, FEMPTY1, FEMPTY2, FEMPTY3, FEMPTY4;
input	[5:0]   FLADJ;
output  EOF1, EOF2, SOFGEN;
output	[13:0]  FRNUM;
output  [10:0]  SOFV;
input   [1:0]   FRLSTSIZE;
input	RUN;			// RUN bit in USBCMD
input	HCHALT;			// HCHALT bit in USBSTS
input	[19:0]	FLBASE;		// periodic frame list base
output	[31:0]	HCIADR1, HCIADR2, HCIADD1, HCIADD2;	// EHCI address, data
output	CMDSTART;		// start MAC cycles
input	MAC_EOT, TXSOF;
output	BUI_GO1, BUI_GO2, BUI_GO3, BUI_GO4, EOT1, EOT2, EOT3, EOT4;
input	TDMAEND1, TDMAEND2, TDMAEND3, TDMAEND4, /*TXTHRESH,*/ CRCERR, BABBLE;
output	RXERR1, RXERR2, RXERR3, RXERR4, HCIMWR1, HCIMWR2;
input	[10:0]	ACTLEN, MAXLEN;
input	/*BOUNDRY,*/ PIDERR, TMOUT, RXNAK, RXNYET, RXSTALL, RXACK;
input	RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXPIDERR;
input	[7:0]	RXPID;
input	[31:0]	WPR1, WPR2;
output	[31:0]  ASYNCLISTADDR;
output	RECLAMATION;
input	TOGMATCH, SPD;
output	ASYNC_ACT, PERIOD_ACT, RUN_C, ROLLOVER_S;
input	WR_ASYNCADDR;
output	[104:0]	TRAN_CMD1, TRAN_CMD2, TRAN_CMD3, TRAN_CMD4;
output	[3:0]	PCIDMA_SEL;//, USBDMA_SEL;
output	[4:0]	USBDMA_SEL;
input	CREQ1, CREQ2, CREQ3, CREQ4;
input	[7:0]	INTTHRESHOLD;	// interrupt threshold
input	USBINT, ERRINT, USBINT_EN, ERRINT_EN;
output	USBINT_S, ERRINT_S;//, IOCSPDINT, USBERRINT;
input   INTASYNC_EN;            // interrupt on async enable
input   INTDOORBELL;            // interrupt on async advance doorbell
input   INTASYNC;               // interrupt on async status
output  INTASYNC_S;             // set interrupt on async status
output  ASYNCINT;               // interrupt on async
output	EHCIEXE;		// EHCI control start processing TDs
input	TEST_PACKET;		// Test_Packet test mode enable
//input	FIFO_OK;		// FIFO control read pipe ready
input	TESTPKTOK;		// Test_Packet FIFO control read pipe ready
input	SWDBG;			// software debug mode
output	HSERR_S;
input	SLAVEMODE;		// select slave mode
output	SLAVE_ACT;		// slave mode is activated
//input	[31:0]	SLQUEUEADDR;	// command queue address
output	BMUCRST_;		// in test modes, reset HS_BMUC
output	[7:0]	SLADDR;		// address for reading command queue
output	SLREAD;			// read sram
input	[31:0]	MDO;
input	DATARDY;		// access command queue ready
output	[31:0]	PERIOD_CMD, ASYNC_CMD;	// commands in slave mode
input	SL_PERIOD;		// execute periodic command in slave mode
input	SL_DATA_PIDERR, SL_ET_ERR, SL_SE_ERR, SL_ACK_ERR;
output	SL_PCIERR;		// PCI error in slave mode
output	SLAVE_ERR;		// error occurs in slave mode
output	[7:0]	SL_ERROFFSET;	// error command address offset in slave mode
//output	EXEITD;			// iTD needs to check DATA PID sequence
output	EHCI_IDLE, TD_IDLE1, TD_IDLE2, TD_IDLE3, TD_IDLE4;
output	TD_PARSE_GO1, TD_PARSE_GO2, TD_PARSE_GO3, TD_PARSE_GO4;
input	[10:0]	RXBCNT;		// RX byte count
input   EN_DBG_PORT;            // DEBUG_PORT enable
input   [31:0]  DBGPORT_SC;     // control/status registers
input   [31:0]  DBGPORT_PID;    // USB PIDs registers
input   [31:0]  DBGPORT_ADDR;   // device address registers
output  DBG_COMPL;              // transaction complete
output  DBG_XACTERR;            // transaction error
output  [7:0]   DBG_RXPID;      // DEBUG_PORT RX PID
output  [3:0]   DBG_RXBCNT;     // DEBUG_PORT RX byte count
output	[51:0]	DBG_TRAN_CMD;	// DEBUG_PORT transaction commands
output	DBG_SEL, EHCI_DBG_MAC_EOT;
input	ATPG_ENI;		// ATPG enable

wire [5:0] FLADJ;
wire [13:0]  FRNUM, FRNUM_AD;
wire [10:0]  SOFV;
wire [31:0]  ADI, ADI1, ADI2;
wire [1:0]   FRLSTSIZE;
wire [3:0] DWCNT;
wire [31:0] HCIADR1, HCIADR2, HCIADD1, HCIADD2;
//wire [31:0] WPR;
//wire [3:0] PCIDMA_SEL, USBDMA_SEL;

//wire GEN_PERR1=1'b0;
//wire PERIOD_ACT=1'b0;

    //sor2b DNT_PERR ( .A(GEN_PERR1), .B(GEN_PERR2), .Y(HSERR_S) );

// split ADI to ADI1 and ADI2
zckbufb DNTAD01 ( .A(ADI[0]), .Y(ADI1[0]) );
zckbufb DNTAD11 ( .A(ADI[1]), .Y(ADI1[1]) );
zckbufb DNTAD21 ( .A(ADI[2]), .Y(ADI1[2]) );
zckbufb DNTAD31 ( .A(ADI[3]), .Y(ADI1[3]) );
zckbufb DNTAD41 ( .A(ADI[4]), .Y(ADI1[4]) );
zckbufb DNTAD51 ( .A(ADI[5]), .Y(ADI1[5]) );
zckbufb DNTAD61 ( .A(ADI[6]), .Y(ADI1[6]) );
zckbufb DNTAD71 ( .A(ADI[7]), .Y(ADI1[7]) );
zckbufb DNTAD81 ( .A(ADI[8]), .Y(ADI1[8]) );
zckbufb DNTAD91 ( .A(ADI[9]), .Y(ADI1[9]) );
zckbufb DNTAD101 ( .A(ADI[10]), .Y(ADI1[10]) );
zckbufb DNTAD111 ( .A(ADI[11]), .Y(ADI1[11]) );
zckbufb DNTAD121 ( .A(ADI[12]), .Y(ADI1[12]) );
zckbufb DNTAD131 ( .A(ADI[13]), .Y(ADI1[13]) );
zckbufb DNTAD141 ( .A(ADI[14]), .Y(ADI1[14]) );
zckbufb DNTAD151 ( .A(ADI[15]), .Y(ADI1[15]) );
zckbufb DNTAD161 ( .A(ADI[16]), .Y(ADI1[16]) );
zckbufb DNTAD171 ( .A(ADI[17]), .Y(ADI1[17]) );
zckbufb DNTAD181 ( .A(ADI[18]), .Y(ADI1[18]) );
zckbufb DNTAD191 ( .A(ADI[19]), .Y(ADI1[19]) );
zckbufb DNTAD201 ( .A(ADI[20]), .Y(ADI1[20]) );
zckbufb DNTAD211 ( .A(ADI[21]), .Y(ADI1[21]) );
zckbufb DNTAD221 ( .A(ADI[22]), .Y(ADI1[22]) );
zckbufb DNTAD231 ( .A(ADI[23]), .Y(ADI1[23]) );
zckbufb DNTAD241 ( .A(ADI[24]), .Y(ADI1[24]) );
zckbufb DNTAD251 ( .A(ADI[25]), .Y(ADI1[25]) );
zckbufb DNTAD261 ( .A(ADI[26]), .Y(ADI1[26]) );
zckbufb DNTAD271 ( .A(ADI[27]), .Y(ADI1[27]) );
zckbufb DNTAD281 ( .A(ADI[28]), .Y(ADI1[28]) );
zckbufb DNTAD291 ( .A(ADI[29]), .Y(ADI1[29]) );
zckbufb DNTAD301 ( .A(ADI[30]), .Y(ADI1[30]) );
zckbufb DNTAD311 ( .A(ADI[31]), .Y(ADI1[31]) );

zckbufb DNTAD02 ( .A(ADI[0]), .Y(ADI2[0]) );
zckbufb DNTAD12 ( .A(ADI[1]), .Y(ADI2[1]) );
zckbufb DNTAD22 ( .A(ADI[2]), .Y(ADI2[2]) );
zckbufb DNTAD32 ( .A(ADI[3]), .Y(ADI2[3]) );
zckbufb DNTAD42 ( .A(ADI[4]), .Y(ADI2[4]) );
zckbufb DNTAD52 ( .A(ADI[5]), .Y(ADI2[5]) );
zckbufb DNTAD62 ( .A(ADI[6]), .Y(ADI2[6]) );
zckbufb DNTAD72 ( .A(ADI[7]), .Y(ADI2[7]) );
zckbufb DNTAD82 ( .A(ADI[8]), .Y(ADI2[8]) );
zckbufb DNTAD92 ( .A(ADI[9]), .Y(ADI2[9]) );
zckbufb DNTAD102 ( .A(ADI[10]), .Y(ADI2[10]) );
zckbufb DNTAD112 ( .A(ADI[11]), .Y(ADI2[11]) );
zckbufb DNTAD122 ( .A(ADI[12]), .Y(ADI2[12]) );
zckbufb DNTAD132 ( .A(ADI[13]), .Y(ADI2[13]) );
zckbufb DNTAD142 ( .A(ADI[14]), .Y(ADI2[14]) );
zckbufb DNTAD152 ( .A(ADI[15]), .Y(ADI2[15]) );
zckbufb DNTAD162 ( .A(ADI[16]), .Y(ADI2[16]) );
zckbufb DNTAD172 ( .A(ADI[17]), .Y(ADI2[17]) );
zckbufb DNTAD182 ( .A(ADI[18]), .Y(ADI2[18]) );
zckbufb DNTAD192 ( .A(ADI[19]), .Y(ADI2[19]) );
zckbufb DNTAD202 ( .A(ADI[20]), .Y(ADI2[20]) );
zckbufb DNTAD212 ( .A(ADI[21]), .Y(ADI2[21]) );
zckbufb DNTAD222 ( .A(ADI[22]), .Y(ADI2[22]) );
zckbufb DNTAD232 ( .A(ADI[23]), .Y(ADI2[23]) );
zckbufb DNTAD242 ( .A(ADI[24]), .Y(ADI2[24]) );
zckbufb DNTAD252 ( .A(ADI[25]), .Y(ADI2[25]) );
zckbufb DNTAD262 ( .A(ADI[26]), .Y(ADI2[26]) );
zckbufb DNTAD272 ( .A(ADI[27]), .Y(ADI2[27]) );
zckbufb DNTAD282 ( .A(ADI[28]), .Y(ADI2[28]) );
zckbufb DNTAD292 ( .A(ADI[29]), .Y(ADI2[29]) );
zckbufb DNTAD302 ( .A(ADI[30]), .Y(ADI2[30]) );
zckbufb DNTAD312 ( .A(ADI[31]), .Y(ADI2[31]) );

    zckbufb DNT_DBG_SEL ( .A(USBDMA_SEL[4]), .Y(DBG_SEL) );

    HS_FMTIMER HS_FMTIMER ( .CLK60M(CLK60M), .TRST_(TRST_), .FLADJ(FLADJ),
	//.REDUCE(REDUCE), .EOF1(EOF1), .EOF2(EOF2), .PRESOF(PRESOF),
	.REDUCE(REDUCE), .EOF1(EHCI_EOF1), .EOF2(EOF2), .PRESOF(PRESOF),
	.FRNUM_PCLK(FRNUM), .PCICLK(EHCIFLOW_PCLK),
	.MAXLEN(MAXLEN), .SOFV(SOFV),
	//.ADI(ADI1), .WR_FRNUM(WR_FRNUM), .RUN(RUN), .HCHALT(HCHALT),
	.ADI(SADI), .WR_FRNUM(WR_FRNUM), .RUN(RUN), .HCHALT(HCHALT),
	.ASYNC_ACT(ASYNC_ACT), .FRNUM_PCLK_LATCH(FRNUM_PCLK_LATCH),
	//.FRLSTSIZE(FRLSTSIZE), .SOFGEN(SOFGEN), .EHCISLEEP(EHCISLEEP),
	.FRLSTSIZE(FRLSTSIZE), .SOFGEN(EHCI_SOFGEN), .EHCISLEEP(EHCISLEEP),
	.EHCIRESTART(EHCIRESTART), .START_EVENT(START_EVENT),
	.FROZEN(FROZEN), .ROLLOVER_S(ROLLOVER_S),
	.INTTHRESHOLD(INTTHRESHOLD), .ITDIOCINT1(ITDIOCINT1),
	.ITDIOCINT2(ITDIOCINT2), .SITDIOCINT1(SITDIOCINT1),
	.SITDIOCINT2(SITDIOCINT2), .USBINT(USBINT),
	/*.IOCSPDINT(IOCSPDINT),*/ .GEN_PERR(HSERR_S), .QHIOCINT1(QHIOCINT1),
	.QHIOCINT2(QHIOCINT2), .QHIOCINT3(QHIOCINT3), .QHIOCINT4(QHIOCINT4),
	.QHERRINT1(QHERRINT1), .QHERRINT2(QHERRINT2), .QHERRINT3(QHERRINT3),
	.QHERRINT4(QHERRINT4), /*.USBERRINT(USBERRINT),*/
	.ERRINT(ERRINT), .INTASYNC(INTASYNC), .ASYNCINT(ASYNCINT),
	.QHASYNCINT(QHASYNCINT), .SWDBG(SWDBG), .MAC_EOT(MAC_EOT),
	.EHCI_MAC_EOT(EHCI_MAC_EOT), .EHCI_DBG_MAC_EOT(EHCI_DBG_MAC_EOT),
	.HSERR_S(HSERR_S),
	.PRESOF_EVAL(PRESOF_EVAL), .HCI_PRESOF(HCI_PRESOF),
	.FRNUM_AD(FRNUM_AD), .LTINT_PCLK(LTINT_PCLK),
	.CMDSTART(CMDSTART), .TXSOF(TXSOF),
	.SLEEPTIME_SEL(SLEEPTIME_SEL), .ATPG_ENI(ATPG_ENI) );

    EHCI_MUX EHCI_MUX ( .GEN_PERR1(GEN_PERR_PER), .GEN_PERR2(GEN_PERR_ASYNC),
	.GEN_PERR(HSERR_S), .RUN_C1(RUN_C1), .RUN_C2(RUN_C2),
	.RUN_C(RUN_C), .FROZEN1(FROZEN1), .FROZEN2(FROZEN2),
	.FROZEN(FROZEN), .ATPG_ENI(ATPG_ENI), .TEST_PACKET(TEST_PACKET),
	.SLAVE_ACT(SLAVE_ACT), .TRST_(TRST_), .BMUCRST_(BMUCRST_),
	.ITDIOCINT_S1(ITDIOCINT_S1), .ITDIOCINT_S2(ITDIOCINT_S2),
	.QHIOCINT_S1(QHIOCINT_S1), .QHIOCINT_S2(QHIOCINT_S2),
	.QHIOCINT_S3(QHIOCINT_S3), .QHIOCINT_S4(QHIOCINT_S4),
	.SITDIOCINT_S1(SITDIOCINT_S1), .SITDIOCINT_S2(SITDIOCINT_S2),
	.ITDERRINT_S1(ITDERRINT_S1), .ITDERRINT_S2(ITDERRINT_S2),
	.QHERRINT_S1(QHERRINT_S1), .QHERRINT_S2(QHERRINT_S2),
	.QHERRINT_S3(QHERRINT_S3), .QHERRINT_S4(QHERRINT_S4),
	.SITDERRINT_S1(SITDERRINT_S1), .SITDERRINT_S2(SITDERRINT_S2),
	.USBINT_S(USBINT_S), .ERRINT_S(ERRINT_S),
	.PER_BUI_GO1(PER_BUI_GO1), .TBUI_GO(TBUI_GO),
	.SLBUI_GO(SLBUI_GO), .SLAVEMODE(SLAVEMODE), .BUI_GO1(BUI_GO1),
	.EHCIFLOW_IDLE(EHCIFLOW_IDLE), .PERIOD_END(PERIOD_END),
	.ASYNC_ACT(ASYNC_ACT), .EHCI_IDLE(EHCI_IDLE)
	/*.PER_HCIADR1(PER_HCIADR1), .SLQUEUEADDR(SLQUEUEADDR),
	.HCIADR1(HCIADR1)*/ );

    EHCIFLOW EHCIFLOW ( .PCIDMA_SEL(PCIDMA_SEL), .USBDMA_SEL(USBDMA_SEL),
	.LIST_SEL(LIST_SEL), .ASYNC_EXE1(ASYNC_EXE1), .ASYNC_EXE2(ASYNC_EXE2),
	.PER_EXE1(PER_EXE1), .PER_EXE2(PER_EXE2), .PERIOD_END(PERIOD_END),
	.PER_CMDSTART_REQ1(PER_CMDSTART_REQ1),
	.PER_CMDSTART_REQ2(PER_CMDSTART_REQ2),
	.ASYNC_CMDSTART_REQ1(QCMDSTART_REQ1),
	.ASYNC_CMDSTART_REQ2(QCMDSTART_REQ2),
	.PER_CMDSTART1(PER_CMDSTART1), .PER_CMDSTART2(PER_CMDSTART2),
	.ASYNC_CMDSTART1(QCMDSTART1), .ASYNC_CMDSTART2(QCMDSTART2),
	.TCMDSTART(TCMDSTART), .TEST_PACKET(TEST_PACKET),
	.SLAVEMODE(SLAVEMODE), .SLCMDSTART(SLCMDSTART),
	.CMDSTART(CMDSTART), .EHCI_MAC_EOT(EHCI_MAC_EOT),
	.CREQ1(CREQ1), .CREQ2(CREQ2), .CREQ3(CREQ3), .CREQ4(CREQ4),
	.ASYNC_EN(ASYNC_EN), .PERIOD_EN(PERIOD_EN), .SOFGEN(SOFGEN),
	//.PRESOF(PRESOF), .EOF1(EOF1), .EOF2(EOF2), .FRNUM(FRNUM),
	.PRESOF(EHCI_DBG_PRESOF), .EOF1(EOF1), .EOF2(EOF2), .FRNUM(FRNUM),
	.PRESOF_EVAL(PRESOF_EVAL), .HCI_PRESOF(HCI_PRESOF),
	//.PERIOD_PRESOF(PERIOD_PRESOF), .TXSOF(TXSOF), .RUN(RUN), .SWDBG(SWDBG),
	.PERIOD_PRESOF(PERIOD_PRESOF), .TXSOF(TXSOF), .RUN(EHCI_DBG_RUN), .SWDBG(SWDBG),
	.EHCIFLOW_IDLE(EHCIFLOW_IDLE), .ASYNC_ACT(ASYNC_ACT),
	.DBG_LIST(DBG_LIST), .DBG_CMDSTART_REQ(DBG_CMDSTART_REQ),
	.DBG_CMDSTART(DBG_CMDSTART), .DBG_ACT(DBG_ACT),
	.EN_DBG_PORT(EN_DBG_PORT),
	.CLK60M(CLK60M), .PCICLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    zivc DNT_DBG_IDLE ( .A(DBG_ACT), .Y(DBG_IDLE) );

    PERIODIC_CTL PERIODIC_CTL ( .PCI1WAIT(PCI1WAIT), .HCIMRDY(HCIMRDY1),
	.RDYACK(RDYACK), .HCICOMPL(HCICOMPL1), .MABORTS(MABORTS),
	.TABORTR(TABORTR), .HCIGNT(HCIGNT1), .EHCIREQ(EHCIREQ1),
	/*.PCICLK(PCICLK),*/ .TRST_(TRST_), .PAROPT(PAROPT), .PERRS(PERRS),
	.SERRS(SERRS), .PMSTR(PMSTR1), .MADDR(MADDR1), .PERIOD_EN(PERIOD_EN),
	.EOFTERM(EOFTERM), .TDMAEND1(TDMAEND1), .TDMAEND2(TDMAEND2),
	.FEMPTY1(FEMPTY1), .FEMPTY2(FEMPTY2), .ADI(ADI2),
	.WPR1(WPR1), .WPR2(WPR2),
	.FLBASE(FLBASE), .FRNUM_AD(FRNUM_AD), .PERIOD_END(PERIOD_END),
	.RUN(RUN), .HCIADR(HCIADR1), .GEN_PERR_PER(GEN_PERR_PER),
	.GEN_PERR(HSERR_S),
	.PER_CMDSTART_REQ1(PER_CMDSTART_REQ1),
	.PER_CMDSTART_REQ2(PER_CMDSTART_REQ2),
	.PER_CMDSTART1(PER_CMDSTART1), .PER_CMDSTART2(PER_CMDSTART2),
	.EHCI_MAC_EOT(EHCI_MAC_EOT), .HCI_PRESOF(PERIOD_PRESOF),
	.BUI_GO1(PER_BUI_GO1), .BUI_GO2(BUI_GO2),
	.TRAN_CMD1(TRAN_CMD1), .TRAN_CMD2(TRAN_CMD2),
	.PER_EXE1(PER_EXE1), .PER_EXE2(PER_EXE2),
	.EOT1(EOT1), .EOT2(EOT2), .RXERR1(RXERR1), .RXERR2(RXERR2),
	.CRCERR(CRCERR), .ACTLEN(ACTLEN), .BABBLE(BABBLE),
	.PIDERR(PIDERR), .TMOUT(TMOUT), .RXNAK(RXNAK), .RXNYET(RXNYET),
	.RXSTALL(RXSTALL), .RXACK(RXACK), .RXDATA0(RXDATA0),
	.RXDATA1(RXDATA1), .RXDATA2(RXDATA2), .RXMDATA(RXMDATA),
	.RXPIDERR(RXPIDERR), .TOGMATCH(TOGMATCH), .SPD(SPD), .RXPID(RXPID),
	.HCIADD(HCIADD1), .HCIMWR(HCIMWR1),
	.PERIOD_ACT(PERIOD_ACT), .RUN_C(RUN_C1),
	.LIST_SEL(LIST_SEL), .USBDMA_SEL(USBDMA_SEL),
	.LTINT_PCLK(LTINT_PCLK),
	.USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN), .USBINT(USBINT),
	.ERRINT(ERRINT), 
	.ITDIOCINT_S1(ITDIOCINT_S1), .ITDIOCINT_S2(ITDIOCINT_S2),
	.ITDERRINT_S1(ITDERRINT_S1), .ITDERRINT_S2(ITDERRINT_S2),
	.QHIOCINT_S1(QHIOCINT_S1), .QHIOCINT_S2(QHIOCINT_S2),
	.QHERRINT_S1(QHERRINT_S1), .QHERRINT_S2(QHERRINT_S2),
	.SITDIOCINT_S1(SITDIOCINT_S1), .SITDIOCINT_S2(SITDIOCINT_S2),
	.SITDERRINT_S1(SITDERRINT_S1), .SITDERRINT_S2(SITDERRINT_S2),
	.ITDIOCINT1(ITDIOCINT1), .ITDIOCINT2(ITDIOCINT2),
	.QHIOCINT1(QHIOCINT1), .QHIOCINT2(QHIOCINT2),
	.SITDIOCINT1(SITDIOCINT1), .SITDIOCINT2(SITDIOCINT2),
	.QHERRINT1(QHERRINT1), .QHERRINT2(QHERRINT2), .FROZEN(FROZEN1),
	//.EHCI_IDLE(EHCI_IDLE), .TDIDLE1(TD_IDLE1), .TDIDLE2(TD_IDLE2),
	.EHCIFLOW_IDLE(EHCIFLOW_IDLE), .TDIDLE1(TD_IDLE1), .TDIDLE2(TD_IDLE2),
	.TD_PARSE_GO1(TD_PARSE_GO1), .TD_PARSE_GO2(TD_PARSE_GO2),
	.SWDBG(SWDBG), .ATPG_ENI(ATPG_ENI),
	.EHCIFLOW_PCLK(EHCIFLOW_PCLK), .EHCI_DMA1_PCLK(EHCI_DMA1_PCLK),
	.EHCI_DMA2_PCLK(EHCI_DMA2_PCLK),
	.EHCIFLOW_CACHE_PCLK(EHCIFLOW_CACHE_PCLK),
	.EHCI_DMA1_CACHE_PCLK(EHCI_DMA1_CACHE_PCLK),
	.EHCI_DMA2_CACHE_PCLK(EHCI_DMA2_CACHE_PCLK),
	.UGNTI_(UGNTI1_), .FRLSTSIZE(FRLSTSIZE) );

    ASYNC_CTL ASYNC_CTL ( .PCI1WAIT(PCI1WAIT), .HCIMRDY(HCIMRDY2),
	.RDYACK(RDYACK), .HCICOMPL(HCICOMPL2), .MABORTS(MABORTS),
	.TABORTR(TABORTR), .HCIGNT(HCIGNT2), .EHCIREQ(EHCIREQ2),
	/*.PCICLK(PCICLK),*/ .TRST_(TRST_), .PAROPT(PAROPT), .PERRS(PERRS),
	.SERRS(SERRS), .PMSTR(PMSTR3), .MADDR(MADDR3), .ASYNC_EN(ASYNC_EN),
	.EOFTERM(EOFTERM), .TDMAEND1(TDMAEND3), .TDMAEND2(TDMAEND4),
	.FEMPTY1(FEMPTY3), .FEMPTY2(FEMPTY4), .ADI(ADI1), .SADI(SADI),
	.RUN(RUN), .HCIADR(HCIADR2), .GEN_PERR_ASYNC(GEN_PERR_ASYNC),
	.GEN_PERR(HSERR_S),
	.QCMDSTART_REQ1(QCMDSTART_REQ1), .QCMDSTART_REQ2(QCMDSTART_REQ2),
	.QCMDSTART1(QCMDSTART1), .QCMDSTART2(QCMDSTART2),
	.EHCI_MAC_EOT(EHCI_MAC_EOT),
	.BUI_GO1(BUI_GO3), .BUI_GO2(BUI_GO4),
	.TRAN_CMD1(TRAN_CMD3), .TRAN_CMD2(TRAN_CMD4),
	.ASYNC_EXE1(ASYNC_EXE1), .ASYNC_EXE2(ASYNC_EXE2),
	.QEOT1(EOT3), .QEOT2(EOT4), .QRXERR1(RXERR3), .QRXERR2(RXERR4),
	.CRCERR(CRCERR), .ACTLEN(ACTLEN), .BABBLE(BABBLE),
	.PIDERR(PIDERR), .TMOUT(TMOUT), .RXNAK(RXNAK), .RXNYET(RXNYET),
	.RXSTALL(RXSTALL), .RXACK(RXACK), .RXDATA0(RXDATA0),
	.RXDATA1(RXDATA1), .RXDATA2(RXDATA2), .RXMDATA(RXMDATA),
	.RXPIDERR(RXPIDERR), .TOGMATCH(TOGMATCH), .SPD(SPD),
	.HCIADD(HCIADD2), .HCIMWR(HCIMWR2), .ASYNCLISTADDR(ASYNCLISTADDR),
	.ASYNC_ACT(ASYNC_ACT), .RUN_C(RUN_C2), .WR_ASYNCADDR(WR_ASYNCADDR),
	.LIST_SEL(LIST_SEL), .RECLAMATION(RECLAMATION),
	.EHCISLEEP(EHCISLEEP), .EHCIRESTART(EHCIRESTART),
	.START_EVENT(START_EVENT), .USBDMA_SEL(USBDMA_SEL),
	.INTASYNC_EN(INTASYNC_EN), .INTASYNC(INTASYNC),
	.INTDOORBELL(INTDOORBELL), .LTINT_PCLK(LTINT_PCLK),
	.INTASYNC_S(INTASYNC_S), .QHASYNCINT(QHASYNCINT),
	.USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN), .USBINT(USBINT),
	.ERRINT(ERRINT), .QHIOCINT_S1(QHIOCINT_S3), .QHIOCINT_S2(QHIOCINT_S4),
	.QHERRINT_S1(QHERRINT_S3), .QHERRINT_S2(QHERRINT_S4),
	.QHIOCINT1(QHIOCINT3), .QHIOCINT2(QHIOCINT4),
	.QHERRINT1(QHERRINT3), .QHERRINT2(QHERRINT4), .FROZEN(FROZEN2),
	.QHIDLE1(TD_IDLE3), .QHIDLE2(TD_IDLE4),
	.QH_PARSE_GO1(TD_PARSE_GO3), .QH_PARSE_GO2(TD_PARSE_GO4),
	.SWDBG(SWDBG), .ATPG_ENI(ATPG_ENI),
	.EHCIFLOW_PCLK(EHCIFLOW_PCLK), .EHCI_DMA1_PCLK(EHCI_DMA3_PCLK),
        .EHCI_DMA2_PCLK(EHCI_DMA4_PCLK),
	.EHCI_DMA1_CACHE_PCLK(EHCI_DMA3_CACHE_PCLK),
        .EHCI_DMA2_CACHE_PCLK(EHCI_DMA4_CACHE_PCLK),
	.UGNTI_(UGNTI3_) );

    DBGCTL DBGCTL ( .EN_DBG_PORT(EN_DBG_PORT),
	.GEN_PERR(HSERR_S), .DBGPORT_SC(DBGPORT_SC),
	.DBGPORT_PID(DBGPORT_PID), .DBGPORT_ADDR(DBGPORT_ADDR),
        .DBG_COMPL(DBG_COMPL), .DBG_XACTERR(DBG_XACTERR),
	.DBG_RXPID(DBG_RXPID), .DBG_RXBCNT(DBG_RXBCNT),
        .DBG_CMDSTART_REQ(DBG_CMDSTART_REQ), .TRAN_CMD(DBG_TRAN_CMD),
	.DBG_ACT(DBG_ACT), .DBG_CMDSTART(DBG_CMDSTART),
        .EHCI_MAC_EOT(EHCI_MAC_EOT), .CRCERR(CRCERR),
	.BABBLE(BABBLE), .PIDERR(PIDERR), .TMOUT(TMOUT),
        .RXACK(RXACK), .RXPID(RXPID), .RXBCNT(RXBCNT),
        .PCICLK(DBG_PCLK), .TRST_(TRST_) );

    DBG_FMTIMER DBG_FMTIMER ( .EN_DBG_PORT(EN_DBG_PORT),
	.DBG_OWNER(DBGPORT_SC[30]), .DBG_ENABLE(DBGPORT_SC[28]), .RUN(RUN),
        .DBG_SOFGEN(DBG_SOFGEN), .EHCI_SOFGEN(EHCI_SOFGEN),
	.SOFGEN(SOFGEN), .EHCI_DBG_RUN(EHCI_DBG_RUN),
        .MAC_EOT(MAC_EOT), .EHCI_DBG_MAC_EOT(EHCI_DBG_MAC_EOT),
	.PRESOF(PRESOF), .EHCI_DBG_PRESOF(EHCI_DBG_PRESOF),
	.EHCI_EOF1(EHCI_EOF1), .EOF1(EOF1),
        .CLK60M(CLK60M), .TRST_(TRST_) );

    TESTPKTCTL TESTPKTCTL ( .PCICLK(EHCIFLOW_PCLK), .TRST_(TRST_),
	.TEST_PACKET(TEST_PACKET), .RUN(RUN), .EHCI_MAC_EOT(EHCI_MAC_EOT),
	.TESTPKTOK(TESTPKTOK), .TBUI_GO(TBUI_GO), .TCMDSTART(TCMDSTART) );

    SLAVECTL SLAVECTL ( .PCICLK(EHCIFLOW_PCLK), .TRST_(TRST_),
	.SLAVEMODE(SLAVEMODE), .EHCI_MAC_EOT(EHCI_MAC_EOT),
	.SLBUI_GO(SLBUI_GO), .SLHCIREQ(SLHCIREQ),
	.SLCMDSTART(SLCMDSTART), .SLREAD(SLREAD), .GEN_PERR(HSERR_S),
	.TDMAEND(TDMAEND1), /*.SLMAXLEN(SLMAXLEN), .SLTRAN_GO(SLTRAN_GO),*/
	.SLAVE_ACT(SLAVE_ACT), .SLADDR(SLADDR), .DATARDY(DATARDY),
	.MDO(MDO), .PERIOD_CMD(PERIOD_CMD), .ASYNC_CMD(ASYNC_CMD),
	.SL_PERIOD(SL_PERIOD), .CRCERR(CRCERR), .PIDERR(PIDERR),
	.SL_DATA_PIDERR(SL_DATA_PIDERR), .SL_ET_ERR(SL_ET_ERR),
	.SL_SE_ERR(SL_SE_ERR), .SL_ACK_ERR(SL_ACK_ERR),
	.SL_PCIERR(SL_PCIERR), .SL_ERROFFSET(SL_ERROFFSET),
	.SLAVE_ERR(SLAVE_ERR) );

endmodule

module PERIODIC_CTL ( PCI1WAIT, HCIMRDY, RDYACK, HCICOMPL,
              MABORTS, TABORTR, HCIGNT, /*PCICLK,*/ TRST_,
              PAROPT, PERRS, SERRS, PMSTR, MADDR, ADI, FLBASE, FRNUM_AD,
	      PERIOD_EN, PERIOD_END, EOFTERM, FEMPTY1, FEMPTY2, EHCIREQ,
	      RUN, HCIADR, HCIADD, PER_CMDSTART_REQ1, PER_CMDSTART_REQ2,
	      PER_CMDSTART1, PER_CMDSTART2, EHCI_MAC_EOT,
	      BUI_GO1, BUI_GO2, TDMAEND1, TDMAEND2, //TXTHRESH,
	      CRCERR, RXERR1, RXERR2, ACTLEN, BABBLE, HCIMWR,
	      WPR1, WPR2, PIDERR, PER_EXE1, PER_EXE2,
	      EOT1, EOT2, LIST_SEL, PERIOD_ACT, HCI_PRESOF,
	      TMOUT, RXNAK, RXNYET, RXSTALL,
	      RXACK, RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXPIDERR, RXPID,
	      TOGMATCH, SPD, GEN_PERR_PER, GEN_PERR,
	      TRAN_CMD1, TRAN_CMD2, USBDMA_SEL,
	      RUN_C, USBINT, ERRINT, USBINT_EN, ERRINT_EN, LTINT_PCLK,
	      ITDIOCINT_S1, ITDIOCINT_S2, ITDERRINT_S1, ITDERRINT_S2,
	      QHIOCINT_S1, QHIOCINT_S2, QHERRINT_S1, QHERRINT_S2,
	      SITDIOCINT_S1, SITDIOCINT_S2, SITDERRINT_S1, SITDERRINT_S2,
	      ITDIOCINT1, ITDIOCINT2, QHIOCINT1, QHIOCINT2,
	      SITDIOCINT1, SITDIOCINT2, QHERRINT1, QHERRINT2, FROZEN,
	      EHCIEXE, SWDBG, EHCIFLOW_IDLE, TDIDLE1, TDIDLE2,
	      TD_PARSE_GO1, TD_PARSE_GO2, ATPG_ENI,
	      EHCIFLOW_PCLK, EHCI_DMA1_PCLK, EHCI_DMA2_PCLK,
	      EHCIFLOW_CACHE_PCLK, EHCI_DMA1_CACHE_PCLK, EHCI_DMA2_CACHE_PCLK,
	      UGNTI_, FRLSTSIZE
            );
input	EHCIFLOW_PCLK, EHCI_DMA1_PCLK, EHCI_DMA2_PCLK;
input	EHCIFLOW_CACHE_PCLK, EHCI_DMA1_CACHE_PCLK, EHCI_DMA2_CACHE_PCLK;
input   PCI1WAIT, RDYACK, MABORTS, TABORTR, PAROPT, PERRS, SERRS, PMSTR;//, MADDR;
output  HCICOMPL, HCIMRDY;
input   /*PCICLK,*/ TRST_, HCIGNT;
input	[31:0]	ADI;		// data bus to latch data
input	[19:0]	FLBASE;		// periodic frame list base
input	[13:0]	FRNUM_AD;
input	PERIOD_EN, EOFTERM, HCI_PRESOF;
output	PERIOD_END, EHCIREQ, GEN_PERR_PER;
input	GEN_PERR, FEMPTY1, FEMPTY2;
input	RUN;			// RUN bit in USBCMD
output	[31:0]	HCIADR, HCIADD;	// EHCI address, data
output	PER_CMDSTART_REQ1, PER_CMDSTART_REQ2;		// start MAC cycles
input	PER_CMDSTART1, PER_CMDSTART2;
input	EHCI_MAC_EOT;
output	BUI_GO1, BUI_GO2;
input	TDMAEND1, TDMAEND2, /*TXTHRESH,*/ CRCERR, BABBLE;
output	RXERR1, RXERR2, HCIMWR;
input	[10:0]	ACTLEN;
output	PER_EXE1, PER_EXE2, EOT1, EOT2;
input	PIDERR, TMOUT, RXNAK, RXNYET, RXSTALL, RXACK;
input	RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXPIDERR;
input	[7:0]	RXPID;
input	[31:0]	WPR1, WPR2;
input	TOGMATCH, SPD, LIST_SEL;
output	PERIOD_ACT, RUN_C;
output	[104:0]	TRAN_CMD1, TRAN_CMD2;
input	[4:0]	USBDMA_SEL;
input	USBINT, ERRINT, USBINT_EN, ERRINT_EN;
output	ITDIOCINT_S1, ITDIOCINT_S2, QHIOCINT_S1, QHIOCINT_S2,
	SITDIOCINT_S1, SITDIOCINT_S2,
	ITDERRINT_S1, ITDERRINT_S2, QHERRINT_S1, QHERRINT_S2,
	SITDERRINT_S1, SITDERRINT_S2, ITDIOCINT1, ITDIOCINT2,
	QHIOCINT1, QHIOCINT2, SITDIOCINT1, SITDIOCINT2,
	QHERRINT1, QHERRINT2;
input	LTINT_PCLK, EHCIFLOW_IDLE;
output	FROZEN;
output	EHCIEXE;		// EHCI control start processing TDs
//input	FIFO_OK;		// FIFO control read pipe ready
input	SWDBG;			// software debug mode
//output	EXEITD;			// iTD needs to check DATA PID sequence
output	TDIDLE1, TDIDLE2;
output	TD_PARSE_GO1, TD_PARSE_GO2;
input	UGNTI_;
output	MADDR;
input	[1:0]	FRLSTSIZE;
input	ATPG_ENI;		// ATPG enable

wire [31:0]  ADI;
wire [3:0] DWCNT;
wire [31:0] DW1_0, DW1_1, DW1_2, DW1_3, DW1_4, DW1_5, DW1_6, DW1_7,
	    DW1_8, DW1_9, DW1_10, DW1_11, DW1_12, DW1_13, DW1_14, DW1_15;
wire [31:0] DW2_0, DW2_1, DW2_2, DW2_3, DW2_4, DW2_5, DW2_6, DW2_7,
	    DW2_8, DW2_9, DW2_10, DW2_11, DW2_12, DW2_13, DW2_14, DW2_15;
wire [31:0] PHCI_DW0, PHCI_DW1;
wire [31:0] IHCIADR1, IHCIADD1, IHCIADR2, IHCIADD2;
wire [31:0] QHCIADR1, QHCIADD1, QHCIADR2, QHCIADD2;
wire [31:0] SIHCIADR1, SIHCIADD1, SIHCIADR2, SIHCIADD2;
wire [3:0] DWNUM, EDWNUM, QHDWNUM1, QHDWNUM2, IDWNUM1, IDWNUM2,
	   SIDWNUM1, SIDWNUM2;
wire [31:0] BUFPTR, /*WPR,*/ IBUFPTR1, IBUFPTR2, INXTLINKPTR;
wire [31:0] UP_DW1_3, UP_DW1_4, UP_DW1_5, UP_DW1_6, UP_DW1_7,
	    UP_DW1_8, UP_DW1_9;
wire [31:0] UP_DW2_3, UP_DW2_4, UP_DW2_5, UP_DW2_6, UP_DW2_7,
	    UP_DW2_8, UP_DW2_9;
wire [31:0] QUP_DW1_3, QUP_DW2_3, SIUP_DW1_3, SIUP_DW2_3;
wire [26:0] CACHE_ADDR1, CACHE_ADDR2;
wire [1:0] NAKCNTSM, NAKCNTSMNXT;
wire [10:0] ACTLEN, ACTLEN1, ACTLEN2;
wire [13:0] FRNUM_PER;
wire [31:0] PERHCIADR;
wire [15:0]  LDW;
wire [3:0] DWOFFSET, QDWOFFSET1, QDWOFFSET2, IDWOFFSET1, IDWOFFSET2,
	   SIDWOFFSET1, SIDWOFFSET2, EDWOFFSET;
wire [104:0] ITRAN_CMD1, ITRAN_CMD2, QTRAN_CMD1, QTRAN_CMD2,
	     SITRAN_CMD1, SITRAN_CMD2;

zckbufb DNTPERR1 ( .A(GEN_PERR), .Y(GEN_PERR_BUF1) );
zckbufb DNTPERR2 ( .A(GEN_PERR), .Y(GEN_PERR_BUF2) );

    HS_PCICTL HS_PCICTL ( .LDW(LDW), .PCI1WAIT(PCI1WAIT), .HCIMRDY(HCIMRDY),
	.RDYACK(RDYACK), .HCICOMPL(HCICOMPL), .PCIEND(PCIEND),
	.MABORTS(MABORTS), .TABORTR(TABORTR), .GEN_PERR(GEN_PERR_PER),
	.HCIGNT(HCIGNT), .PCICLK(EHCIFLOW_PCLK), .TRST_(TRST_), .PAROPT(PAROPT),
	.PERRS(PERRS), .SERRS(SERRS), .PMSTR(PMSTR), //.MADDR(MADDR), 
	.EDWNUM(EDWNUM), .DWCNT(DWCNT), .HCIMWR(HCIMWR),
	.EDWOFFSET(EDWOFFSET), .ATPG_ENI(ATPG_ENI),
	.MADDR(MADDR), .UGNTI_(UGNTI_) );

    //sivb DNT_CACHEN1 ( .A(CACHE_SEL), .Y(CACHE_EN1) );
    //sycbufb DNT_CACHEN2 ( .A(CACHE_SEL), .Y(CACHE_EN2) );

    PHCI_CACHE PHCI_CACHE ( .LDW(LDW), .ADI(ADI),
	.PCICLK(EHCIFLOW_CACHE_PCLK),
	.TRST_(TRST_), .DW0(PHCI_DW0), .DW1(PHCI_DW1),
	.CACHE_EN(PCACHE_EN), .ATPG_ENI(ATPG_ENI) );

    PERIODIC_CACHE PERIODIC_CACHE1 ( .LDW(LDW), .ADI(ADI),
	.PCICLK(EHCI_DMA1_CACHE_PCLK), .TRST_(TRST_), .DW0(DW1_0), .DW1(DW1_1),
	.DW2(DW1_2), .DW3(DW1_3), .DW4(DW1_4), .DW5(DW1_5),
	.DW6(DW1_6), .DW7(DW1_7), .DW8(DW1_8), .DW9(DW1_9),
	.DW10(DW1_10), .DW11(DW1_11), .DW12(DW1_12), .DW13(DW1_13),
	.DW14(DW1_14), .DW15(DW1_15),
	.CACHEPHASE(CACHEPHASE1),
	.UP_DW3(UP_DW1_3), .UP_DW4(UP_DW1_4), .UP_DW5(UP_DW1_5),
	.UP_DW6(UP_DW1_6), .UP_DW7(UP_DW1_7), .UP_DW8(UP_DW1_8),
	.UP_DW9(UP_DW1_9), .UP_LDW3(UP_LDW1_3),
	.UP_LDW4(UP_LDW1_4), .UP_LDW5(UP_LDW1_5),
	.UP_LDW6(UP_LDW1_6), .UP_LDW7(UP_LDW1_7),
	.UP_LDW8(UP_LDW1_8), .UP_LDW9(UP_LDW1_9),
	.CACHE_EN(CACHE_EN1), .ATPG_ENI(ATPG_ENI) );

    PERIODIC_CACHE PERIODIC_CACHE2 ( .LDW(LDW), .ADI(ADI),
        .PCICLK(EHCI_DMA2_CACHE_PCLK), .TRST_(TRST_), .DW0(DW2_0), .DW1(DW2_1),
	.DW2(DW2_2), .DW3(DW2_3), .DW4(DW2_4), .DW5(DW2_5),
	.DW6(DW2_6), .DW7(DW2_7), .DW8(DW2_8), .DW9(DW2_9),
	.DW10(DW2_10), .DW11(DW2_11), .DW12(DW2_12), .DW13(DW2_13),
	.DW14(DW2_14), .DW15(DW2_15),
        .CACHEPHASE(CACHEPHASE2),
        .UP_DW3(UP_DW2_3), .UP_DW4(UP_DW2_4), .UP_DW5(UP_DW2_5),
	.UP_DW6(UP_DW2_6), .UP_DW7(UP_DW2_7), .UP_DW8(UP_DW2_8),
	.UP_DW9(UP_DW2_9), .UP_LDW3(UP_LDW2_3),
	.UP_LDW4(UP_LDW2_4), .UP_LDW5(UP_LDW2_5),
	.UP_LDW6(UP_LDW2_6), .UP_LDW7(UP_LDW2_7),
	.UP_LDW8(UP_LDW2_8), .UP_LDW9(UP_LDW2_9),
        .CACHE_EN(CACHE_EN2), .ATPG_ENI(ATPG_ENI) );

    PERIODICFLOW PERIODICFLOW ( .PERIOD_EN(PERIOD_EN), .PCIEND(PCIEND),
	.GEN_PERR(GEN_PERR_BUF1), .PERIOD_END(PERIOD_END),
	.HCI_PRESOF(HCI_PRESOF), .PHCI_PRESOF(PHCI_PRESOF), 
	.RUN(RUN), .DWNUM(DWNUM),  .PERIOD_ACT(PERIOD_ACT),
	.EHCIREQ(EHCIREQ), .PARSETDEND1(PARSETDEND1),
	.PARSETDEND2(PARSETDEND2), .TDPARSING1(TDPARSING1),
	.TDPARSING2(TDPARSING2), .EXEITD1(EXEITD1), .EXEITD2(EXEITD2),
	.EXEQH1(EXEQH1), .EXEQH2(EXEQH2), .EXESITD1(EXESITD1), 
	.EXESITD2(EXESITD2), .ITDIDLE1(ITDIDLE1), .ITDIDLE2(ITDIDLE2),
	.QHIDLE1(QHIDLE1), .QHIDLE2(QHIDLE2), .SITDIDLE1(SITDIDLE1),
	.SITDIDLE2(SITDIDLE2), .TDIDLE1(TDIDLE1), .TDIDLE2(TDIDLE2),
	.PHCI_DW0(PHCI_DW0), .PHCI_DW1(PHCI_DW1),
	.DW1_0(DW1_0), .DW2_0(DW2_0),
	.CACHE_INVALID1(CACHE_INVALID1), .CACHE_INVALID2(CACHE_INVALID2),
	.TD_CACHE_EN1(TD_CACHE_EN1), .TD_CACHE_EN2(TD_CACHE_EN2),
	.TD_PARSE_GO1(TD_PARSE_GO1), .TD_PARSE_GO2(TD_PARSE_GO2),
	.DWOFFSET(DWOFFSET), .PCACHE_EN(PCACHE_EN),
	.CACHE_EN1(CACHE_EN1), .CACHE_EN2(CACHE_EN2),
	.TD_ACT1(TD_ACT1), .TD_ACT2(TD_ACT2),
	.PER_EXE1(PER_EXE1), .PER_EXE2(PER_EXE2),
	.TDHCIREQ1(TDHCIREQ1), .TDHCIREQ2(TDHCIREQ2),
	.TDHCIGNT1(TDHCIGNT1), .TDHCIGNT2(TDHCIGNT2),
	.CACHE_ADDR1(CACHE_ADDR1), .CACHE_ADDR2(CACHE_ADDR2),
	.TDEXE1(TDEXE1), .TDEXE2(TDEXE2), .PERHCIADR(PERHCIADR),
	.FRNUM(FRNUM_AD), .FRNUM_PER(FRNUM_PER), .FLBASE(FLBASE),
	.LIST_SEL(LIST_SEL), .LTINT_PCLK(LTINT_PCLK),
	.SWDBG(SWDBG), .RUN_C(RUN_C), .FROZEN(FROZEN),
	.TDCMDSTART1(PER_CMDSTART1), .TDCMDSTART2(PER_CMDSTART2),
	//.RECOVERYMODE(RECOVERYMODE), .EHCI_IDLE(EHCI_IDLE),
	.RECOVERYMODE(RECOVERYMODE), .EHCIFLOW_IDLE(EHCIFLOW_IDLE),
	.PCICLK(EHCIFLOW_PCLK), .TRST_(TRST_), .FRLSTSIZE(FRLSTSIZE) );

    ITDCTL ITDCTL1 ( .ITD_PARSE_GO(ITD_PARSE_GO1), .PARSEITDEND(PARSEITDEND1),
	.ITDPARSING(ITDPARSING1), .ITDIDLE(ITDIDLE1), .FRNUM(FRNUM_PER),
	.DW0(DW1_0), .DW1(DW1_1), .DW2(DW1_2), .DW3(DW1_3), .DW4(DW1_4),
	.DW5(DW1_5), .DW6(DW1_6), .DW7(DW1_7), .DW8(DW1_8), .DW9(DW1_9),
	.DW10(DW1_10), .DW11(DW1_11), .DW12(DW1_12), .DW13(DW1_13),
	.DW14(DW1_14), .DW15(DW1_15), .GEN_PERR(GEN_PERR_BUF1),
	.PCIEND(IPCIEND1), .IHCIREQ(IHCIREQ1), .IDWNUM(IDWNUM1),
	.IDWOFFSET(IDWOFFSET1), .IHCIADR(IHCIADR1), .IHCIADD(IHCIADD1),
	.IHCIMWR(IHCIMWR1), .TRAN_CMD(ITRAN_CMD1), .ITD_ACT(ITD_ACT1),
	.IBUI_GO(IBUI_GO1), .CACHE_ADDR(CACHE_ADDR1),
	.CACHE_INVALID(ICACHE_INVALID1), .WPR(WPR1),
	.CRCERR(CRCERR1), .ACTLEN(ACTLEN1), .BABBLE(BABBLE1),
	.PIDERR(PIDERR1), .TMOUT(TMOUT1), .RXDATA0(RXDATA01),
	.RXDATA1(RXDATA11), .RXDATA2(RXDATA21), .RXPID(RXPID),
	.TOGMATCH(TOGMATCH1), .SPD(SPD1), .EHCI_MAC_EOT(ITD_MAC_EOT1),
	.FEMPTY(FEMPTY1), .TDMAEND(TDMAEND1), .IRXERR(IRXERR1),
	.ICMDSTART_REQ(ICMDSTART_REQ1), .ICMDSTART(ICMDSTART1),
	.IEOT(IEOT1), .HCI_PRESOF(HCI_PRESOF), .LTINT_PCLK(LTINT_PCLK),
	.USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN),
	.USBINT(USBINT), .ERRINT(ERRINT),
	.ITDIOCINT_S(ITDIOCINT_S1), .ITDERRINT_S(ITDERRINT_S1),
	.ITDIOCINT(ITDIOCINT1), .RECOVERYMODE(RECOVERYMODE),
	.PCICLK(EHCI_DMA1_PCLK), .EHCIFLOW_PCLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    ITDCTL ITDCTL2 ( .ITD_PARSE_GO(ITD_PARSE_GO2), .PARSEITDEND(PARSEITDEND2),
	.ITDPARSING(ITDPARSING2), .ITDIDLE(ITDIDLE2), .FRNUM(FRNUM_PER),
	.DW0(DW2_0), .DW1(DW2_1), .DW2(DW2_2), .DW3(DW2_3), .DW4(DW2_4),
	.DW5(DW2_5), .DW6(DW2_6), .DW7(DW2_7), .DW8(DW2_8), .DW9(DW2_9),
	.DW10(DW2_10), .DW11(DW2_11), .DW12(DW2_12), .DW13(DW2_13),
	.DW14(DW2_14), .DW15(DW2_15), .GEN_PERR(GEN_PERR_BUF2),
	.PCIEND(IPCIEND2), .IHCIREQ(IHCIREQ2), .IDWNUM(IDWNUM2),
	.IDWOFFSET(IDWOFFSET2), .IHCIADR(IHCIADR2), .IHCIADD(IHCIADD2),
	.IHCIMWR(IHCIMWR2), .TRAN_CMD(ITRAN_CMD2), .ITD_ACT(ITD_ACT2),
	.IBUI_GO(IBUI_GO2), .CACHE_ADDR(CACHE_ADDR2),
	.CACHE_INVALID(ICACHE_INVALID2), .WPR(WPR2),
	.CRCERR(CRCERR2), .ACTLEN(ACTLEN2), .BABBLE(BABBLE2),
	.PIDERR(PIDERR2), .TMOUT(TMOUT2), .RXDATA0(RXDATA02),
	.RXDATA1(RXDATA12), .RXDATA2(RXDATA22), .RXPID(RXPID),
	.TOGMATCH(TOGMATCH2), .SPD(SPD2), .EHCI_MAC_EOT(ITD_MAC_EOT2),
	.FEMPTY(FEMPTY2), .TDMAEND(TDMAEND2), .IRXERR(IRXERR2),
	.ICMDSTART_REQ(ICMDSTART_REQ2), .ICMDSTART(ICMDSTART2),
	.IEOT(IEOT2), .HCI_PRESOF(HCI_PRESOF), .LTINT_PCLK(LTINT_PCLK),
	.USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN),
	.USBINT(USBINT), .ERRINT(ERRINT),
	.ITDIOCINT_S(ITDIOCINT_S2), .ITDERRINT_S(ITDERRINT_S2),
	.ITDIOCINT(ITDIOCINT2), .RECOVERYMODE(RECOVERYMODE),
	.PCICLK(EHCI_DMA2_PCLK), .EHCIFLOW_PCLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    PQHCTL PQHCTL1 ( .QH_PARSE_GO(QH_PARSE_GO1), .QHPARSING(QHPARSING1),
	.PARSEQHEND(PARSEQHEND1), .DW0(DW1_0), .DW1(DW1_1), .DW2(DW1_2),
	.DW3(DW1_3), .DW4(DW1_4), .DW5(DW1_5), .DW6(DW1_6), .DW7(DW1_7),
	.DW8(DW1_8), .DW9(DW1_9), .DW10(DW1_10), .DW11(DW1_11),
	.GEN_PERR(GEN_PERR_BUF1), .PCIEND(QPCIEND1), .DWCNT(DWCNT),
	.UP_DW3(QUP_DW1_3), .UP_DW6(UP_DW1_6),
	.UP_DW7(UP_DW1_7), .UP_DW8(UP_DW1_8), .UP_DW9(UP_DW1_9),
	.UP_LDW3(QUP_LDW1_3), .UP_LDW6(UP_LDW1_6),
	.UP_LDW7(UP_LDW1_7), .UP_LDW8(UP_LDW1_8), .UP_LDW9(UP_LDW1_9),
	.CACHE_INVALID(QCACHE_INVALID1), .FRNUM(FRNUM_PER),
	.QHCIMWR(QHCIMWR1), .QHIDLE(QHIDLE1),
	.QHCIREQ(QHCIREQ1), .QHDWNUM(QHDWNUM1), .QDWOFFSET(QDWOFFSET1),
	.TRAN_CMD(QTRAN_CMD1), .QHCIADR(QHCIADR1), .QHCIADD(QHCIADD1),
	.CACHEPHASE(QCACHEPHASE1), .QBUI_GO(QBUI_GO1), .QH_ACT(QH_ACT1),
	.CRCERR(CRCERR1), .ACTLEN(ACTLEN1), .BABBLE(BABBLE1),
        .PIDERR(PIDERR1), .TMOUT(TMOUT1), .RXNAK(RXNAK1), .RXNYET(RXNYET1),
        .RXSTALL(RXSTALL1), .RXACK(RXACK1), .RXDATA0(RXDATA01),
        .RXDATA1(RXDATA11), .RXMDATA(RXMDATA1), .RXPIDERR(RXPIDERR1),
	.TOGMATCH(TOGMATCH1), .SPD(SPD1),
	.FEMPTY(FEMPTY1), .EHCI_MAC_EOT(QH_MAC_EOT1),
	.QCMDSTART_REQ(QCMDSTART_REQ1), .QCMDSTART(QCMDSTART1),
	.TDMAEND(TDMAEND1), .QEOT(QEOT1), .QRXERR(QRXERR1),
	.CACHE_ADDR(CACHE_ADDR1), .QTDEXE(QTDEXE1), .HCI_PRESOF(PHCI_PRESOF),
	.LTINT_PCLK(LTINT_PCLK), .USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN),
	.USBINT(USBINT), .ERRINT(ERRINT), .QHIOCINT_S(QHIOCINT_S1),
	.QHERRINT_S(QHERRINT_S1), .QHIOCINT(QHIOCINT1), .QHERRINT(QHERRINT1),
	.RECOVERYMODE(RECOVERYMODE), .PCICLK(EHCI_DMA1_PCLK),
	.EHCIFLOW_PCLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    PQHCTL PQHCTL2 ( .QH_PARSE_GO(QH_PARSE_GO2), .QHPARSING(QHPARSING2),
	.PARSEQHEND(PARSEQHEND2), .DW0(DW2_0), .DW1(DW2_1), .DW2(DW2_2),
	.DW3(DW2_3), .DW4(DW2_4), .DW5(DW2_5), .DW6(DW2_6), .DW7(DW2_7),
	.DW8(DW2_8), .DW9(DW2_9), .DW10(DW2_10), .DW11(DW2_11),
	.GEN_PERR(GEN_PERR_BUF2), .PCIEND(QPCIEND2), .DWCNT(DWCNT),
	.UP_DW3(QUP_DW2_3), .UP_DW6(UP_DW2_6),
	.UP_DW7(UP_DW2_7), .UP_DW8(UP_DW2_8), .UP_DW9(UP_DW2_9),
	.UP_LDW3(QUP_LDW2_3), .UP_LDW6(UP_LDW2_6),
	.UP_LDW7(UP_LDW2_7), .UP_LDW8(UP_LDW2_8), .UP_LDW9(UP_LDW2_9),
	.CACHE_INVALID(QCACHE_INVALID2), .FRNUM(FRNUM_PER),
	.QHCIMWR(QHCIMWR2), .QHIDLE(QHIDLE2),
	.QHCIREQ(QHCIREQ2), .QHDWNUM(QHDWNUM2), .QDWOFFSET(QDWOFFSET2),
	.TRAN_CMD(QTRAN_CMD2), .QHCIADR(QHCIADR2), .QHCIADD(QHCIADD2),
	.CACHEPHASE(QCACHEPHASE2), .QBUI_GO(QBUI_GO2), .QH_ACT(QH_ACT2),
	.CRCERR(CRCERR2), .ACTLEN(ACTLEN2), .BABBLE(BABBLE2),
        .PIDERR(PIDERR2), .TMOUT(TMOUT2), .RXNAK(RXNAK2), .RXNYET(RXNYET2),
        .RXSTALL(RXSTALL2), .RXACK(RXACK2), .RXDATA0(RXDATA02),
        .RXDATA1(RXDATA12), .RXMDATA(RXMDATA2), .RXPIDERR(RXPIDERR2),
	.TOGMATCH(TOGMATCH2), .SPD(SPD2),
	.FEMPTY(FEMPTY2), .EHCI_MAC_EOT(QH_MAC_EOT2),
	.QCMDSTART_REQ(QCMDSTART_REQ2), .QCMDSTART(QCMDSTART2),
	.TDMAEND(TDMAEND2), .QEOT(QEOT2), .QRXERR(QRXERR2),
	.CACHE_ADDR(CACHE_ADDR2), .QTDEXE(QTDEXE2), .HCI_PRESOF(PHCI_PRESOF),
	.LTINT_PCLK(LTINT_PCLK), .USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN),
	.USBINT(USBINT), .ERRINT(ERRINT), .QHIOCINT_S(QHIOCINT_S2),
	.QHERRINT_S(QHERRINT_S2), .QHIOCINT(QHIOCINT2), .QHERRINT(QHERRINT2),
	.RECOVERYMODE(RECOVERYMODE), .PCICLK(EHCI_DMA2_PCLK),
	.EHCIFLOW_PCLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    SITDCTL SITDCTL1 ( .SITD_PARSE_GO(SITD_PARSE_GO1),
	.PARSESITDEND(PARSESITDEND1), .SITDPARSING(SITDPARSING1),
	.SITDIDLE(SITDIDLE1), .FRNUM(FRNUM_PER), .DWCNT(DWCNT),
	.DW0(DW1_0), .DW1(DW1_1), .DW2(DW1_2), .DW3(DW1_3), .DW4(DW1_4),
	.DW5(DW1_5), .DW6(DW1_6), .DW7(DW1_7), .DW8(DW1_8), .DW9(DW1_9),
	.DW10(DW1_10), .DW11(DW1_11), .DW12(DW1_12), .DW13(DW1_13),
	.GEN_PERR(GEN_PERR_BUF1), .UP_DW3(SIUP_DW1_3), .UP_DW4(UP_DW1_4),
	.UP_DW5(UP_DW1_5), .UP_LDW3(SIUP_LDW1_3), .UP_LDW4(UP_LDW1_4),
	.UP_LDW5(UP_LDW1_5), .CACHEPHASE(SICACHEPHASE1),
	.CACHE_INVALID(SICACHE_INVALID1),
	.PCIEND(SIPCIEND1), .SIHCIREQ(SIHCIREQ1), .SIDWNUM(SIDWNUM1),
	.SIDWOFFSET(SIDWOFFSET1), .SIHCIADR(SIHCIADR1), .SIHCIADD(SIHCIADD1),
	.SIHCIMWR(SIHCIMWR1), .TRAN_CMD(SITRAN_CMD1), .SITD_ACT(SITD_ACT1),
	.SIBUI_GO(SIBUI_GO1), .CACHE_ADDR(CACHE_ADDR1),
	.CRCERR(CRCERR1), .ACTLEN(ACTLEN1), .BABBLE(BABBLE1),
	.PIDERR(PIDERR1), .TMOUT(TMOUT1), .RXDATA0(RXDATA01),
	.RXDATA1(RXDATA11), .RXMDATA(RXMDATA1), .RXNYET(RXNYET1),
	.RXPIDERR(RXPIDERR1), .EHCI_MAC_EOT(SITD_MAC_EOT1),
	.FEMPTY(FEMPTY1), .TDMAEND(TDMAEND1), .SIRXERR(SIRXERR1),
	.SICMDSTART_REQ(SICMDSTART_REQ1), .SICMDSTART(SICMDSTART1),
	.SIEOT(SIEOT1), .HCI_PRESOF(HCI_PRESOF), .LTINT_PCLK(LTINT_PCLK),
	.USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN),
	.USBINT(USBINT), .ERRINT(ERRINT),
	.SITDIOCINT_S(SITDIOCINT_S1), .SITDERRINT_S(SITDERRINT_S1),
	.SITDIOCINT(SITDIOCINT1), .RECOVERYMODE(RECOVERYMODE),
	.PCICLK(EHCI_DMA1_PCLK), .EHCIFLOW_PCLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    SITDCTL SITDCTL2 ( .SITD_PARSE_GO(SITD_PARSE_GO2),
	.PARSESITDEND(PARSESITDEND2), .SITDPARSING(SITDPARSING2),
	.SITDIDLE(SITDIDLE2), .FRNUM(FRNUM_PER), .DWCNT(DWCNT),
	.DW0(DW2_0), .DW1(DW2_1), .DW2(DW2_2), .DW3(DW2_3), .DW4(DW2_4),
	.DW5(DW2_5), .DW6(DW2_6), .DW7(DW2_7), .DW8(DW2_8), .DW9(DW2_9),
	.DW10(DW2_10), .DW11(DW2_11), .DW12(DW2_12), .DW13(DW2_13),
	.GEN_PERR(GEN_PERR_BUF2), .UP_DW3(SIUP_DW2_3), .UP_DW4(UP_DW2_4),
	.UP_DW5(UP_DW2_5), .UP_LDW3(SIUP_LDW2_3), .UP_LDW4(UP_LDW2_4),
	.UP_LDW5(UP_LDW2_5), .CACHEPHASE(SICACHEPHASE2),
	.CACHE_INVALID(SICACHE_INVALID2),
	.PCIEND(SIPCIEND2), .SIHCIREQ(SIHCIREQ2), .SIDWNUM(SIDWNUM2),
	.SIDWOFFSET(SIDWOFFSET2), .SIHCIADR(SIHCIADR2), .SIHCIADD(SIHCIADD2),
	.SIHCIMWR(SIHCIMWR2), .TRAN_CMD(SITRAN_CMD2), .SITD_ACT(SITD_ACT2),
	.SIBUI_GO(SIBUI_GO2), .CACHE_ADDR(CACHE_ADDR2),
	.CRCERR(CRCERR2), .ACTLEN(ACTLEN2), .BABBLE(BABBLE2),
	.PIDERR(PIDERR2), .TMOUT(TMOUT2), .RXDATA0(RXDATA02),
	.RXDATA1(RXDATA12), .RXMDATA(RXMDATA2), .RXNYET(RXNYET2),
	.RXPIDERR(RXPIDERR2), .EHCI_MAC_EOT(SITD_MAC_EOT2),
	.FEMPTY(FEMPTY2), .TDMAEND(TDMAEND2), .SIRXERR(SIRXERR2),
	.SICMDSTART_REQ(SICMDSTART_REQ2), .SICMDSTART(SICMDSTART2),
	.SIEOT(SIEOT2), .HCI_PRESOF(HCI_PRESOF), .LTINT_PCLK(LTINT_PCLK),
	.USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN),
	.USBINT(USBINT), .ERRINT(ERRINT),
	.SITDIOCINT_S(SITDIOCINT_S2), .SITDERRINT_S(SITDERRINT_S2),
	.SITDIOCINT(SITDIOCINT2), .RECOVERYMODE(RECOVERYMODE),
	.PCICLK(EHCI_DMA2_PCLK), .EHCIFLOW_PCLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    PERIODIC_ADCTL PERIODIC_ADCTL ( .PCICLK(EHCIFLOW_PCLK), .TRST_(TRST_),
	.DWCNT(DWCNT), .RUN(RUN), .ADI(ADI), .PERHCIADR(PERHCIADR),
	//.FLBASE(FLBASE),
	//.FRNUM_AD(FRNUM_PER),
	//.DW1_0(DW1_0), .DW2_0(DW2_0),
	//.PARSEQHEND1(PARSEQHEND1), .PARSEQHEND2(PARSEQHEND2),
	.EXEITD1(EXEITD1), .EXEITD2(EXEITD2),
	.EXESITD1(EXESITD1), .EXESITD2(EXESITD2),
	.TDHCIGNT1(TDHCIGNT1), .TDHCIGNT2(TDHCIGNT2),
	.IHCIADR1(IHCIADR1), .IHCIADR2(IHCIADR2),
	.QHCIADR1(QHCIADR1), .QHCIADR2(QHCIADR2),
	.SIHCIADR1(SIHCIADR1), .SIHCIADR2(SIHCIADR2),
	.HCIADR(HCIADR),
	.IHCIADD1(IHCIADD1), .IHCIADD2(IHCIADD2),
	.QHCIADD1(QHCIADD1), .QHCIADD2(QHCIADD2),
	.SIHCIADD1(SIHCIADD1), .SIHCIADD2(SIHCIADD2),
	.HCIADD(HCIADD) );

    PERIODIC_MUX PERIODIC_MUX ( .TD_CACHE_EN1(TD_CACHE_EN1),
	.TD_CACHE_EN2(TD_CACHE_EN2), .EXEITD1(EXEITD1), .EXEITD2(EXEITD2),
	.EXEQH1(EXEQH1), .EXEQH2(EXEQH2), .EXESITD1(EXESITD1),
	.EXESITD2(EXESITD2),
	.DWNUM(DWNUM), .IDWNUM1(IDWNUM1), .QHDWNUM1(QHDWNUM1),
	.SIDWNUM1(SIDWNUM1), .IDWNUM2(IDWNUM2), .QHDWNUM2(QHDWNUM2),
	.SIDWNUM2(SIDWNUM2), .EDWNUM(EDWNUM),
	.DWOFFSET(DWOFFSET),
	.IDWOFFSET1(IDWOFFSET1), .IDWOFFSET2(IDWOFFSET2),
	.QHDWOFFSET1(QDWOFFSET1), .QHDWOFFSET2(QDWOFFSET2),
	.SIDWOFFSET1(SIDWOFFSET1), .SIDWOFFSET2(SIDWOFFSET2),
	.EDWOFFSET(EDWOFFSET), 
	.QUP_DW1_3(QUP_DW1_3), .QUP_DW2_3(QUP_DW2_3),
	.SIUP_DW1_3(SIUP_DW1_3), .SIUP_DW2_3(SIUP_DW2_3),
	.UP_DW1_3(UP_DW1_3), .UP_DW2_3(UP_DW2_3),
	.QUP_LDW1_3(QUP_LDW1_3), .QUP_LDW2_3(QUP_LDW2_3),
	.SIUP_LDW1_3(SIUP_LDW1_3), .SIUP_LDW2_3(SIUP_LDW2_3),
	.UP_LDW1_3(UP_LDW1_3), .UP_LDW2_3(UP_LDW2_3),
	.QCACHEPHASE1(QCACHEPHASE1), .QCACHEPHASE2(QCACHEPHASE2),
	.SICACHEPHASE1(SICACHEPHASE1), .SICACHEPHASE2(SICACHEPHASE2),
	.CACHEPHASE1(CACHEPHASE1), .CACHEPHASE2(CACHEPHASE2),
	.TDHCIREQ1(TDHCIREQ1), .TDHCIREQ2(TDHCIREQ2),
	.IHCIREQ1(IHCIREQ1), .IHCIREQ2(IHCIREQ2), .QHCIREQ1(QHCIREQ1),
	.QHCIREQ2(QHCIREQ2), .SIHCIREQ1(SIHCIREQ1), .SIHCIREQ2(SIHCIREQ2),
	.EHCI_MAC_EOT(EHCI_MAC_EOT),
	.TD_ACT1(TD_ACT1), .TD_ACT2(TD_ACT2), .ITD_ACT1(ITD_ACT1),
	.ITD_ACT2(ITD_ACT2), .QH_ACT1(QH_ACT1), .QH_ACT2(QH_ACT2),
	.SITD_ACT1(SITD_ACT1), .SITD_ACT2(SITD_ACT2),
	.ITD_MAC_EOT1(ITD_MAC_EOT1), .ITD_MAC_EOT2(ITD_MAC_EOT2),
	.QH_MAC_EOT1(QH_MAC_EOT1), .QH_MAC_EOT2(QH_MAC_EOT2),
	.SITD_MAC_EOT1(SITD_MAC_EOT1), .SITD_MAC_EOT2(SITD_MAC_EOT2),
	.TDHCIGNT1(TDHCIGNT1), .TDHCIGNT2(TDHCIGNT2),
	.IMWR1(IHCIMWR1), .IMWR2(IHCIMWR2),
	.SIMWR1(SIHCIMWR1), .SIMWR2(SIHCIMWR2),
	.QHMWR1(QHCIMWR1), .QHMWR2(QHCIMWR2), .HCIMWR(HCIMWR),
	.PARSEITDEND1(PARSEITDEND1), .PARSEITDEND2(PARSEITDEND2),
	.PARSEQHEND1(PARSEQHEND1), .PARSEQHEND2(PARSEQHEND2),
	.PARSESITDEND1(PARSESITDEND1), .PARSESITDEND2(PARSESITDEND2),
	.PARSETDEND1(PARSETDEND1), .PARSETDEND2(PARSETDEND2),
	.ITDPARSING1(ITDPARSING1), .ITDPARSING2(ITDPARSING2),
	.QHPARSING1(QHPARSING1), .QHPARSING2(QHPARSING2),
	.SITDPARSING1(SITDPARSING1), .SITDPARSING2(SITDPARSING2),
	.TDPARSING1(TDPARSING1), .TDPARSING2(TDPARSING2),
	.TD_PARSE_GO1(TD_PARSE_GO1), .TD_PARSE_GO2(TD_PARSE_GO2),
	.ITD_PARSE_GO1(ITD_PARSE_GO1), .ITD_PARSE_GO2(ITD_PARSE_GO2),
	.QH_PARSE_GO1(QH_PARSE_GO1), .QH_PARSE_GO2(QH_PARSE_GO2),
	.SITD_PARSE_GO1(SITD_PARSE_GO1), .SITD_PARSE_GO2(SITD_PARSE_GO2),
	.ICACHE_INVALID1(ICACHE_INVALID1), .ICACHE_INVALID2(ICACHE_INVALID2),
	.QCACHE_INVALID1(QCACHE_INVALID1), .QCACHE_INVALID2(QCACHE_INVALID2),
	.SICACHE_INVALID1(SICACHE_INVALID1),
	.SICACHE_INVALID2(SICACHE_INVALID2),
	.CACHE_INVALID1(CACHE_INVALID1), .CACHE_INVALID2(CACHE_INVALID2),
	.ICMDSTART_REQ1(ICMDSTART_REQ1), .ICMDSTART_REQ2(ICMDSTART_REQ2),
	.QCMDSTART_REQ1(QCMDSTART_REQ1), .QCMDSTART_REQ2(QCMDSTART_REQ2),
	.SICMDSTART_REQ1(SICMDSTART_REQ1), .SICMDSTART_REQ2(SICMDSTART_REQ2),
	.PER_CMDSTART_REQ1(PER_CMDSTART_REQ1),
	.PER_CMDSTART_REQ2(PER_CMDSTART_REQ2),
	.PER_CMDSTART1(PER_CMDSTART1), .PER_CMDSTART2(PER_CMDSTART2),
	.ICMDSTART1(ICMDSTART1), .ICMDSTART2(ICMDSTART2),
	.QCMDSTART1(QCMDSTART1), .QCMDSTART2(QCMDSTART2),
	.SICMDSTART1(SICMDSTART1), .SICMDSTART2(SICMDSTART2),
	.PCIEND(PCIEND), .IPCIEND1(IPCIEND1), .IPCIEND2(IPCIEND2),
	.QPCIEND1(QPCIEND1), .QPCIEND2(QPCIEND2),
	.SIPCIEND1(SIPCIEND1), .SIPCIEND2(SIPCIEND2), .USBDMA_SEL(USBDMA_SEL),
	.ITRAN_CMD1(ITRAN_CMD1), .ITRAN_CMD2(ITRAN_CMD2),
	.QTRAN_CMD1(QTRAN_CMD1), .QTRAN_CMD2(QTRAN_CMD2),
	.SITRAN_CMD1(SITRAN_CMD1), .SITRAN_CMD2(SITRAN_CMD2),
	.TRAN_CMD1(TRAN_CMD1), .TRAN_CMD2(TRAN_CMD2),
	.IBUI_GO1(IBUI_GO1), .IBUI_GO2(IBUI_GO2),
	.QBUI_GO1(QBUI_GO1), .QBUI_GO2(QBUI_GO2),
	.SIBUI_GO1(SIBUI_GO1), .SIBUI_GO2(SIBUI_GO2),
	.BUI_GO1(BUI_GO1), .BUI_GO2(BUI_GO2),
	.IRXERR1(IRXERR1), .IRXERR2(IRXERR2),
	.QRXERR1(QRXERR1), .QRXERR2(QRXERR2),
	.SIRXERR1(SIRXERR1), .SIRXERR2(SIRXERR2),
	.RXERR1(RXERR1), .RXERR2(RXERR2),
	.IEOT1(IEOT1), .IEOT2(IEOT2), .QEOT1(QEOT1), .QEOT2(QEOT2),
	.SIEOT1(SIEOT1), .SIEOT2(SIEOT2), .EOT1(EOT1), .EOT2(EOT2),
	.CRCERR(CRCERR), .BABBLE(BABBLE), .PIDERR(PIDERR), .TMOUT(TMOUT),
	.TOGMATCH(TOGMATCH), .RXNAK(RXNAK), .RXNYET(RXNYET),
	.RXSTALL(RXSTALL), .RXACK(RXACK), .RXDATA0(RXDATA0),
	.RXDATA1(RXDATA1), .RXDATA2(RXDATA2), .RXMDATA(RXMDATA),
	.RXPIDERR(RXPIDERR), .SPD(SPD), .ACTLEN(ACTLEN),
	.CRCERR1(CRCERR1), .BABBLE1(BABBLE1), .PIDERR1(PIDERR1),
	.TMOUT1(TMOUT1), .TOGMATCH1(TOGMATCH1), .RXNAK1(RXNAK1),
	.RXNYET1(RXNYET1), .RXSTALL1(RXSTALL1), .RXACK1(RXACK1),
	.RXDATA01(RXDATA01), .RXDATA11(RXDATA11),
	.RXDATA21(RXDATA21), .RXMDATA1(RXMDATA1),
	.RXPIDERR1(RXPIDERR1), .SPD1(SPD1), .ACTLEN1(ACTLEN1),
	.CRCERR2(CRCERR2), .BABBLE2(BABBLE2), .PIDERR2(PIDERR2),
	.TMOUT2(TMOUT2), .TOGMATCH2(TOGMATCH2), .RXNAK2(RXNAK2),
	.RXNYET2(RXNYET2), .RXSTALL2(RXSTALL2), .RXACK2(RXACK2),
	.RXDATA02(RXDATA02), .RXDATA12(RXDATA12),
	.RXDATA22(RXDATA22), .RXMDATA2(RXMDATA2),
	.RXPIDERR2(RXPIDERR2), .SPD2(SPD2), .ACTLEN2(ACTLEN2) );

endmodule

module ASYNC_CTL ( PCI1WAIT, HCIMRDY, RDYACK, HCICOMPL,
              MABORTS, TABORTR, HCIGNT, /*PCICLK,*/ TRST_,
              PAROPT, PERRS, SERRS, PMSTR, MADDR, ADI, SADI,
	      ASYNC_EN, EOFTERM, FEMPTY1, FEMPTY2, EHCIREQ,
	      RUN, HCIADR, HCIADD, QCMDSTART_REQ1, QCMDSTART_REQ2,
	      QCMDSTART1, QCMDSTART2, EHCI_MAC_EOT,
	      BUI_GO1, BUI_GO2, TDMAEND1, TDMAEND2, //TXTHRESH,
	      CRCERR, QRXERR1, QRXERR2, ACTLEN, BABBLE, HCIMWR,
	      /*BOUNDRY, WPR,*/ PIDERR, ASYNC_EXE1, ASYNC_EXE2,
	      QEOT1, QEOT2, LIST_SEL, EHCISLEEP, EHCIRESTART, START_EVENT,
	      ASYNCLISTADDR, RECLAMATION, TMOUT, RXNAK, RXNYET, RXSTALL,
	      RXACK, RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXPIDERR, RXPID,
	      TOGMATCH, SPD, GEN_PERR_ASYNC, GEN_PERR,
	      TRAN_CMD1, TRAN_CMD2, USBDMA_SEL,
	      ASYNC_ACT, RUN_C, WR_ASYNCADDR,
	      USBINT, ERRINT,
	      USBINT_EN, ERRINT_EN, INTDOORBELL, INTASYNC_EN,
	      INTASYNC_S, INTASYNC, LTINT_PCLK, QHASYNCINT,
	      QHIOCINT_S1, QHIOCINT_S2, QHERRINT_S1, QHERRINT_S2,
	      QHIOCINT1, QHIOCINT2, QHERRINT1, QHERRINT2, FROZEN,
	      EHCIEXE, SWDBG, QHIDLE1, QHIDLE2, QH_PARSE_GO1, QH_PARSE_GO2,
	      EHCIFLOW_PCLK, EHCI_DMA1_PCLK, EHCI_DMA2_PCLK,
	      EHCI_DMA1_CACHE_PCLK, EHCI_DMA2_CACHE_PCLK,
	      UGNTI_, ATPG_ENI
            );
input	EHCIFLOW_PCLK, EHCI_DMA1_PCLK, EHCI_DMA2_PCLK;
input	EHCI_DMA1_CACHE_PCLK, EHCI_DMA2_CACHE_PCLK;
input   PCI1WAIT, RDYACK, MABORTS, TABORTR, PAROPT, PERRS, SERRS, PMSTR;//, MADDR;
output  HCICOMPL, HCIMRDY;
input   /*PCICLK,*/ TRST_, HCIGNT;
input	[31:0]	ADI;		// data bus to latch data
input	[31:0]	SADI;		// data bus to latch data
input	ASYNC_EN, EOFTERM;
output	EHCIREQ, GEN_PERR_ASYNC;
input	GEN_PERR, FEMPTY1, FEMPTY2;
input	RUN;			// RUN bit in USBCMD
output	[31:0]	HCIADR, HCIADD;	// EHCI address, data
output	QCMDSTART_REQ1, QCMDSTART_REQ2;		// start MAC cycles
input	QCMDSTART1, QCMDSTART2;
input	EHCI_MAC_EOT;
output	BUI_GO1, BUI_GO2;
input	TDMAEND1, TDMAEND2, /*TXTHRESH,*/ CRCERR, BABBLE;
output	QRXERR1, QRXERR2, HCIMWR;
input	[10:0]	ACTLEN;
output	ASYNC_EXE1, ASYNC_EXE2, QEOT1, QEOT2;
input	/*BOUNDRY,*/ PIDERR, TMOUT, RXNAK, RXNYET, RXSTALL, RXACK;
input	RXDATA0, RXDATA1, RXDATA2, RXMDATA, RXPIDERR;
input	[7:0]	RXPID;
//input	[31:0]	WPR;
output	[31:0]  ASYNCLISTADDR;
output	RECLAMATION, EHCISLEEP, START_EVENT;
input	TOGMATCH, SPD, LIST_SEL, EHCIRESTART;
output	ASYNC_ACT, RUN_C;
input	WR_ASYNCADDR;
output	[104:0]	TRAN_CMD1, TRAN_CMD2;
input	[4:0]	USBDMA_SEL;
input	USBINT, ERRINT, USBINT_EN, ERRINT_EN;
output	QHIOCINT_S1, QHIOCINT_S2, QHERRINT_S1, QHERRINT_S2,
	QHIOCINT1, QHIOCINT2, QHERRINT1, QHERRINT2;
input   INTASYNC_EN;            // interrupt on async enable
input   INTDOORBELL;            // interrupt on async advance doorbell
input   INTASYNC;               // interrupt on async status
output  INTASYNC_S;             // set interrupt on async status
output  QHASYNCINT;             // interrupt on async
input	LTINT_PCLK;
output	FROZEN;
output	EHCIEXE;		// EHCI control start processing TDs
//input	FIFO_OK;		// FIFO control read pipe ready
input	SWDBG;			// software debug mode
output	QHIDLE1, QHIDLE2;
output	QH_PARSE_GO1, QH_PARSE_GO2;
input	UGNTI_;
output	MADDR;
input	ATPG_ENI;		// ATPG enable

wire [31:0]  ADI;
wire [3:0] DWCNT;
wire [31:0] DW1_0, DW1_1, DW1_2, DW1_3, DW1_4, DW1_5, DW1_6,
	    DW1_7, DW1_8, DW1_9, DW1_10, DW1_11;
wire [31:0] DW2_0, DW2_1, DW2_2, DW2_3, DW2_4, DW2_5, DW2_6,
	    DW2_7, DW2_8, DW2_9, DW2_10, DW2_11;
wire [31:0] QHCIADR1, QHCIADD1, QHCIADR2, QHCIADD2;
wire [3:0] DWNUM, EDWNUM, QHDWNUM1, QHDWNUM2;
wire [31:0] BUFPTR, /*WPR,*/ IBUFPTR1, IBUFPTR2, INXTLINKPTR;
wire [31:0] UP_DW1_3, UP_DW1_5, UP_DW1_6, UP_DW1_7;
wire [31:0] UP_DW2_3, UP_DW2_5, UP_DW2_6, UP_DW2_7;
wire [26:0] CACHE_ADDR1, CACHE_ADDR2;
wire [1:0] NAKCNTSM, NAKCNTSMNXT;
wire [10:0] ACTLEN, ACTLEN1, ACTLEN2;

wire [15:0]  LDW;
wire [3:0] DWOFFSET, QDWOFFSET1, QDWOFFSET2, EDWOFFSET;
//wire HCIMWR=1'b0;
//wire PARK_EN = 1'b0;
//wire [1:0] PARKCNT=2'b0;

zckbufb DNTPERR ( .A(GEN_PERR), .Y(GEN_PERR_BUF) );

    HS_PCICTL HS_PCICTL ( .LDW(LDW), .PCI1WAIT(PCI1WAIT), .HCIMRDY(HCIMRDY),
	.RDYACK(RDYACK), .HCICOMPL(HCICOMPL), .PCIEND(PCIEND),
	.MABORTS(MABORTS), .TABORTR(TABORTR), .GEN_PERR(GEN_PERR_ASYNC),
	.HCIGNT(HCIGNT), .PCICLK(EHCIFLOW_PCLK), .TRST_(TRST_), .PAROPT(PAROPT),
	.PERRS(PERRS), .SERRS(SERRS), .PMSTR(PMSTR), //.MADDR(MADDR), 
	.EDWNUM(EDWNUM), .DWCNT(DWCNT), .HCIMWR(HCIMWR),
	.EDWOFFSET(EDWOFFSET), .ATPG_ENI(ATPG_ENI),
	.MADDR(MADDR), .UGNTI_(UGNTI_) );

    zivb DNT_CACHEN1 ( .A(CACHE_SEL), .Y(CACHE_EN1) );
    zckbufb DNT_CACHEN2 ( .A(CACHE_SEL), .Y(CACHE_EN2) );

    ASYNC_CACHE ASYNC_CACHE1 ( .LDW(LDW), .ADI(ADI),
	.PCICLK(EHCI_DMA1_CACHE_PCLK), .TRST_(TRST_), .DW0(DW1_0), .DW1(DW1_1),
	.DW2(DW1_2), .DW3(DW1_3), .DW4(DW1_4), .DW5(DW1_5),
	.DW6(DW1_6), .DW7(DW1_7), .DW8(DW1_8), .DW9(DW1_9),
	.DW10(DW1_10), .DW11(DW1_11),
	.CACHEPHASE(CACHEPHASE1),
	.UP_DW3(UP_DW1_3), .UP_DW5(UP_DW1_5), .UP_DW6(UP_DW1_6),
	.UP_DW7(UP_DW1_7), .UP_LDW3(UP_LDW1_3), .UP_LDW5(UP_LDW1_5),
	.UP_LDW6(UP_LDW1_6), .UP_LDW7(UP_LDW1_7),
	.CACHE_EN(CACHE_EN1), .ATPG_ENI(ATPG_ENI) );

    ASYNC_CACHE ASYNC_CACHE2 ( .LDW(LDW), .ADI(ADI),
        .PCICLK(EHCI_DMA2_CACHE_PCLK), .TRST_(TRST_), .DW0(DW2_0), .DW1(DW2_1),
	.DW2(DW2_2), .DW3(DW2_3), .DW4(DW2_4), .DW5(DW2_5),
	.DW6(DW2_6), .DW7(DW2_7), .DW8(DW2_8), .DW9(DW2_9),
	.DW10(DW2_10), .DW11(DW2_11),
        .CACHEPHASE(CACHEPHASE2),
        .UP_DW3(UP_DW2_3), .UP_DW5(UP_DW2_5), .UP_DW6(UP_DW2_6),
	.UP_DW7(UP_DW2_7), .UP_LDW3(UP_LDW2_3), .UP_LDW5(UP_LDW2_5),
	.UP_LDW6(UP_LDW2_6), .UP_LDW7(UP_LDW2_7),
        .CACHE_EN(CACHE_EN2), .ATPG_ENI(ATPG_ENI) );

/*
    ASYC_CACHE_MUX ASYC_CACHE_MUX ( .DW1_0(DW1_0), .DW1_1(DW1_1),
	.DW1_2(DW1_2), .DW1_3(DW1_3), .DW1_4(DW1_4), .DW1_5(DW1_5),
	.DW1_6(DW1_6), .DW1_7(DW1_7), .DW1_8(DW1_8), .DW1_9(DW1_9),
	.DW1_10(DW1_10), .DW1_11(DW1_11),
	.DW2_0(DW2_0), .DW2_1(DW2_1),
        .DW2_2(DW2_2), .DW2_3(DW2_3), .DW2_4(DW2_4), .DW2_5(DW2_5),
        .DW2_6(DW2_6), .DW2_7(DW2_7), .DW2_8(DW2_8), .DW2_9(DW2_9),
        .DW2_10(DW2_10), .DW2_11(DW2_11),
	.DW0(DW0), .DW1(DW1), .DW2(DW2),
	.DW3(DW3), .DW4(DW4), .DW5(DW5), .DW6(DW6), .DW7(DW7), .DW8(DW8),
	.DW9(DW9), .DW10(DW10), .DW11(DW11), .CACHE_SEL(CACHE_SEL) );
*/

    ASYNCFLOW ASYNCFLOW ( .ASYNC_EN(ASYNC_EN), .PCIEND(PCIEND),
	.GEN_PERR(GEN_PERR_BUF), //.HCI_PRESOF(HCI_PRESOF),
	.RUN(RUN), .DWNUM(DWNUM),  .ASYNC_ACT(ASYNC_ACT),
	.EHCIREQ(EHCIREQ), .PARSEQHEND1(PARSEQHEND1),
	.PARSEQHEND2(PARSEQHEND2), .QHPARSING1(QHPARSING1),
	.QHPARSING2(QHPARSING2), .QHIDLE1(QHIDLE1), .QHIDLE2(QHIDLE2),
	.QH_CACHE_EN1(QH_CACHE_EN1), .QH_CACHE_EN2(QH_CACHE_EN2),
	.QH_PARSE_GO1(QH_PARSE_GO1), .QH_PARSE_GO2(QH_PARSE_GO2),
	.DWOFFSET(DWOFFSET), .CACHE_SEL(CACHE_SEL),
	.ASYNCLISTADDR(ASYNCLISTADDR),
	.QH_ACT1(QH_ACT1), .QH_ACT2(QH_ACT2),
	.ASYNC_EXE1(ASYNC_EXE1), .ASYNC_EXE2(ASYNC_EXE2),
	.QHCIREQ1(QHCIREQ1), .QHCIREQ2(QHCIREQ2),
	.QHCIGNT1(QHCIGNT1), .QHCIGNT2(QHCIGNT2),
	.CACHE_ADDR1(CACHE_ADDR1), .CACHE_ADDR2(CACHE_ADDR2),
	.QTDEXE1(QTDEXE1), .QTDEXE2(QTDEXE2),
	.CACHE_INVALID1(CACHE_INVALID1), .CACHE_INVALID2(CACHE_INVALID2),
	.HEADSEEN1(HEADSEEN1), .HEADSEEN2(HEADSEEN2),
	.LIST_SEL(LIST_SEL), .RECLAMATION(RECLAMATION),
	.ASYNC_EMPTY1(ASYNC_EMPTY1), .ASYNC_EMPTY2(ASYNC_EMPTY2),
	.EHCISLEEP(EHCISLEEP), .EHCIRESTART(EHCIRESTART),
	.START_EVENT(START_EVENT),
	.NAKCNTSM(NAKCNTSM), .NAKCNTSMNXT(NAKCNTSMNXT),
	.INTASYNC_EN(INTASYNC_EN), .INTASYNC(INTASYNC),
	.INTDOORBELL(INTDOORBELL), .LTINT_PCLK(LTINT_PCLK),
	.INTASYNC_S(INTASYNC_S), .QHASYNCINT(QHASYNCINT),
	.SWDBG(SWDBG), .RUN_C(RUN_C), .FROZEN(FROZEN),
	.QCMDSTART1(QCMDSTART1), .QCMDSTART2(QCMDSTART2),
	.PCICLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    AQHCTL AQHCTL1 ( .QH_PARSE_GO(QH_PARSE_GO1), .QHPARSING(QHPARSING1),
	.PARSEQHEND(PARSEQHEND1), .DW0(DW1_0), .DW1(DW1_1), .DW2(DW1_2),
	.DW3(DW1_3), .DW4(DW1_4), .DW5(DW1_5), .DW6(DW1_6), .DW7(DW1_7),
	.DW8(DW1_8), .DW9(DW1_9), .DW10(DW1_10), .DW11(DW1_11),
	.GEN_PERR(GEN_PERR_BUF), .PCIEND(QPCIEND1), .DWCNT(DWCNT),
	//.PARK_EN(PARK_EN), .PARKCNT(PARKCNT),
	.UP_DW3(UP_DW1_3), .UP_DW5(UP_DW1_5), .UP_DW6(UP_DW1_6),
	.UP_DW7(UP_DW1_7),
	.UP_LDW3(UP_LDW1_3), .UP_LDW5(UP_LDW1_5), .UP_LDW6(UP_LDW1_6),
	.UP_LDW7(UP_LDW1_7), .CACHE_INVALID(CACHE_INVALID1),
	.QHCIMWR(QHCIMWR1), .QHIDLE(QHIDLE1),
	.QHCIREQ(QHCIREQ1), .QHDWNUM(QHDWNUM1), .QDWOFFSET(QDWOFFSET1),
	.TRAN_CMD(TRAN_CMD1), .QHCIADR(QHCIADR1), .QHCIADD(QHCIADD1),
	.CACHEPHASE(CACHEPHASE1), .QBUI_GO(BUI_GO1), .QH_ACT(QH_ACT1),
	.CRCERR(CRCERR1), .ACTLEN(ACTLEN1), .BABBLE(BABBLE1),
        .PIDERR(PIDERR1), .TMOUT(TMOUT1), .RXNAK(RXNAK1), .RXNYET(RXNYET1),
        .RXSTALL(RXSTALL1), .RXACK(RXACK1), .RXDATA0(RXDATA01),
        .RXDATA1(RXDATA11), .RXPIDERR(RXPIDERR1),
	.TOGMATCH(TOGMATCH1), .SPD(SPD1),
	.FEMPTY(FEMPTY1), .EHCI_MAC_EOT(QH_MAC_EOT1),
	.QCMDSTART_REQ(QCMDSTART_REQ1), .QCMDSTART(QCMDSTART1),
	.TDMAEND(TDMAEND1), .QEOT(QEOT1), .QRXERR(QRXERR1),
	.CACHE_ADDR(CACHE_ADDR1),
	.QTDEXE(QTDEXE1), .HEADSEEN(HEADSEEN1), .RECLAMATION(RECLAMATION),
	.ASYNC_EMPTY(ASYNC_EMPTY1),
	.NAKCNTSM(NAKCNTSM), .NAKCNTSMNXT(NAKCNTSMNXT),
	.LTINT_PCLK(LTINT_PCLK), .USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN),
	.USBINT(USBINT), .ERRINT(ERRINT), .QHIOCINT_S(QHIOCINT_S1),
	.QHERRINT_S(QHERRINT_S1), .QHIOCINT(QHIOCINT1), .QHERRINT(QHERRINT1),
	.PCICLK(EHCI_DMA1_PCLK), .EHCIFLOW_PCLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    AQHCTL AQHCTL2 ( .QH_PARSE_GO(QH_PARSE_GO2), .QHPARSING(QHPARSING2),
	.PARSEQHEND(PARSEQHEND2), .DW0(DW2_0), .DW1(DW2_1), .DW2(DW2_2),
	.DW3(DW2_3), .DW4(DW2_4), .DW5(DW2_5), .DW6(DW2_6), .DW7(DW2_7),
	.DW8(DW2_8), .DW9(DW2_9), .DW10(DW2_10), .DW11(DW2_11),
	.GEN_PERR(GEN_PERR_BUF), .PCIEND(QPCIEND2), .DWCNT(DWCNT),
	//.PARK_EN(PARK_EN), .PARKCNT(PARKCNT),
	.UP_DW3(UP_DW2_3), .UP_DW5(UP_DW2_5), .UP_DW6(UP_DW2_6),
	.UP_DW7(UP_DW2_7),
	.UP_LDW3(UP_LDW2_3), .UP_LDW5(UP_LDW2_5), .UP_LDW6(UP_LDW2_6),
	.UP_LDW7(UP_LDW2_7), .CACHE_INVALID(CACHE_INVALID2),
	.QHCIMWR(QHCIMWR2), .QHIDLE(QHIDLE2),
	.QHCIREQ(QHCIREQ2), .QHDWNUM(QHDWNUM2), .QDWOFFSET(QDWOFFSET2),
	.TRAN_CMD(TRAN_CMD2), .QHCIADR(QHCIADR2), .QHCIADD(QHCIADD2),
	.CACHEPHASE(CACHEPHASE2), .QBUI_GO(BUI_GO2), .QH_ACT(QH_ACT2),
	.CRCERR(CRCERR2), .ACTLEN(ACTLEN2), .BABBLE(BABBLE2),
        .PIDERR(PIDERR2), .TMOUT(TMOUT2), .RXNAK(RXNAK2), .RXNYET(RXNYET2),
        .RXSTALL(RXSTALL2), .RXACK(RXACK2), .RXDATA0(RXDATA02),
        .RXDATA1(RXDATA12), .RXPIDERR(RXPIDERR2),
	.TOGMATCH(TOGMATCH2), .SPD(SPD2),
	.FEMPTY(FEMPTY2), .EHCI_MAC_EOT(QH_MAC_EOT2),
	.QCMDSTART_REQ(QCMDSTART_REQ2), .QCMDSTART(QCMDSTART2),
	.TDMAEND(TDMAEND2), .QEOT(QEOT2), .QRXERR(QRXERR2),
	.CACHE_ADDR(CACHE_ADDR2),
	.QTDEXE(QTDEXE2), .HEADSEEN(HEADSEEN2), .RECLAMATION(RECLAMATION),
	.ASYNC_EMPTY(ASYNC_EMPTY2),
	.NAKCNTSM(NAKCNTSM), .NAKCNTSMNXT(NAKCNTSMNXT),
	.LTINT_PCLK(LTINT_PCLK), .USBINT_EN(USBINT_EN), .ERRINT_EN(ERRINT_EN),
	.USBINT(USBINT), .ERRINT(ERRINT), .QHIOCINT_S(QHIOCINT_S2),
	.QHERRINT_S(QHERRINT_S2), .QHIOCINT(QHIOCINT2), .QHERRINT(QHERRINT2),
	.PCICLK(EHCI_DMA2_PCLK), .EHCIFLOW_PCLK(EHCIFLOW_PCLK), .TRST_(TRST_) );

    ASYNC_ADCTL ASYNC_ADCTL ( .PCICLK(EHCIFLOW_PCLK), .TRST_(TRST_),
	.DWCNT(DWCNT), .WR_ASYNCADDR(WR_ASYNCADDR), .RUN(RUN),
	.ADI(SADI), .ASYNC_ACT(ASYNC_ACT), .ASYNC_EN(ASYNC_EN),
	.ASYNCLISTADDR(ASYNCLISTADDR), .DW1_0(DW1_0), .DW2_0(DW2_0),
	.PARSEQHEND1(PARSEQHEND1), .PARSEQHEND2(PARSEQHEND2),
	.QHCIGNT1(QHCIGNT1), .QHCIGNT2(QHCIGNT2),
	.QHCIADR1(QHCIADR1), .QHCIADR2(QHCIADR2), .HCIADR(HCIADR),
	.QHCIADD1(QHCIADD1), .QHCIADD2(QHCIADD2), .HCIADD(HCIADD),
	.ASYNC_EMPTY1(ASYNC_EMPTY1), .ASYNC_EMPTY2(ASYNC_EMPTY2) );

    ASYNC_MUX ASYNC_MUX ( .QH_CACHE_EN1(QH_CACHE_EN1),
	.QH_CACHE_EN2(QH_CACHE_EN2), .DWNUM(DWNUM),
	.QHDWNUM1(QHDWNUM1), .QHDWNUM2(QHDWNUM2), .EDWNUM(EDWNUM),
	.DWOFFSET(DWOFFSET), .QDWOFFSET1(QDWOFFSET1), .QDWOFFSET2(QDWOFFSET2),
	.EDWOFFSET(EDWOFFSET), /*.HCIREQ(HCIREQ), .QHCIREQ1(QHCIREQ1),
	.QHCIREQ2(QHCIREQ2), .EHCIREQ(EHCIREQ),*/ .EHCI_MAC_EOT(EHCI_MAC_EOT),
	.QH_ACT1(QH_ACT1), .QH_ACT2(QH_ACT2), .QH_MAC_EOT1(QH_MAC_EOT1),
	.QHCIGNT1(QHCIGNT1), .QHCIGNT2(QHCIGNT2),
	.QHCIMWR1(QHCIMWR1), .QHCIMWR2(QHCIMWR2), .HCIMWR(HCIMWR),
	.QH_MAC_EOT2(QH_MAC_EOT2), .PCIEND(PCIEND), .QPCIEND1(QPCIEND1),
	.QPCIEND2(QPCIEND2), .USBDMA_SEL(USBDMA_SEL),
	.CRCERR(CRCERR), .BABBLE(BABBLE), .PIDERR(PIDERR), .TMOUT(TMOUT),
	.TOGMATCH(TOGMATCH), .RXNAK(RXNAK), .RXNYET(RXNYET),
	.RXSTALL(RXSTALL), .RXACK(RXACK), .RXDATA0(RXDATA0),
	.RXDATA1(RXDATA1), .RXPIDERR(RXPIDERR), .SPD(SPD), .ACTLEN(ACTLEN),
	.CRCERR1(CRCERR1), .BABBLE1(BABBLE1), .PIDERR1(PIDERR1),
	.TMOUT1(TMOUT1), .TOGMATCH1(TOGMATCH1), .RXNAK1(RXNAK1),
	.RXNYET1(RXNYET1), .RXSTALL1(RXSTALL1), .RXACK1(RXACK1),
	.RXDATA01(RXDATA01), .RXDATA11(RXDATA11), .RXPIDERR1(RXPIDERR1),
	.SPD1(SPD1), .ACTLEN1(ACTLEN1),
	.CRCERR2(CRCERR2), .BABBLE2(BABBLE2), .PIDERR2(PIDERR2),
	.TMOUT2(TMOUT2), .TOGMATCH2(TOGMATCH2), .RXNAK2(RXNAK2),
	.RXNYET2(RXNYET2), .RXSTALL2(RXSTALL2), .RXACK2(RXACK2),
	.RXDATA02(RXDATA02), .RXDATA12(RXDATA12), .RXPIDERR2(RXPIDERR2),
	.SPD2(SPD2), .ACTLEN2(ACTLEN2) );

endmodule



module HS_INTF ( PSADO31, PSADO30, PSADO29, PSADO28, PSADO27, PSADO26, PSADO25, 
    PSADO24, PSADO23, PSADO22, PSADO21, PSADO20, PSADO19, PSADO18, PSADO17, 
    PSADO16, PSADO15, PSADO14, PSADO13, PSADO12, PSADO11, PSADO10, PSADO9, 
    PSADO8, PSADO7, PSADO6, PSADO5, PSADO4, PSADO3, PSADO2, PSADO1, PSADO0, 
    UHIT, ULRDY, CFGW, REGW, REGR, REGADS, RDYACK, IRDYI_, TRDYI_, AD31I, 
    AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I, AD23I, AD22I, AD21I, 
    AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, AD14I, AD13I, AD12I, AD11I, 
    AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I, LCMD0, 
    REGD31, REGD30, REGD29, REGD28, REGD27, REGD26, REGD25, REGD24, REGD23, 
    REGD22, REGD21, REGD20, REGD19, REGD18, REGD17, REGD16, REGD15, REGD14, 
    REGD13, REGD12, REGD11, REGD10, REGD9, REGD8, REGD7, REGD6, REGD5, REGD4, 
    REGD3, REGD2, REGD1, REGD0, CFGD31, CFGD30, CFGD29, CFGD28, CFGD27, CFGD26, 
    CFGD25, CFGD24, CFGD23, CFGD22, CFGD21, CFGD20, CFGD19, CFGD18, CFGD17, 
    CFGD16, CFGD15, CFGD14, CFGD13, CFGD12, CFGD11, CFGD10, CFGD9, CFGD8, 
    CFGD7, CFGD6, CFGD5, CFGD4, CFGD3, CFGD2, CFGD1, CFGD0, CBE3I_, CBE2I_, 
    CBE1I_, CBE0I_, IOBA31, IOBA30, IOBA29, IOBA28, IOBA27, IOBA26, IOBA25, 
    IOBA24, IOBA23, IOBA22, IOBA21, IOBA20, IOBA19, IOBA18, IOBA17, IOBA16, 
    IOBA15, IOBA14, IOBA13, IOBA12, IOBA11, IOBA10, IOBA9, IOBA8, UADS, 
    IOSPACE, PMSTR, EN_EHCI, HRST_, PCICLK, ADS, ADRG, IDSELI, FUNCSEL, PA7I, 
    PA6I, PA5I, PA4I, PA3I, PA2I );
input  [2:0] FUNCSEL;
input  IRDYI_, TRDYI_, AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I, 
    AD23I, AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, AD14I, 
    AD13I, AD12I, AD11I, AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, 
    AD1I, AD0I, REGD31, REGD30, REGD29, REGD28, REGD27, REGD26, REGD25, REGD24, 
    REGD23, REGD22, REGD21, REGD20, REGD19, REGD18, REGD17, REGD16, REGD15, 
    REGD14, REGD13, REGD12, REGD11, REGD10, REGD9, REGD8, REGD7, REGD6, REGD5, 
    REGD4, REGD3, REGD2, REGD1, REGD0, CFGD31, CFGD30, CFGD29, CFGD28, CFGD27, 
    CFGD26, CFGD25, CFGD24, CFGD23, CFGD22, CFGD21, CFGD20, CFGD19, CFGD18, 
    CFGD17, CFGD16, CFGD15, CFGD14, CFGD13, CFGD12, CFGD11, CFGD10, CFGD9, 
    CFGD8, CFGD7, CFGD6, CFGD5, CFGD4, CFGD3, CFGD2, CFGD1, CFGD0, CBE3I_, 
    CBE2I_, CBE1I_, CBE0I_, IOBA31, IOBA30, IOBA29, IOBA28, IOBA27, IOBA26, 
    IOBA25, IOBA24, IOBA23, IOBA22, IOBA21, IOBA20, IOBA19, IOBA18, IOBA17, 
    IOBA16, IOBA15, IOBA14, IOBA13, IOBA12, IOBA11, IOBA10, IOBA9, IOBA8, UADS, 
    IOSPACE, PMSTR, EN_EHCI, HRST_, PCICLK, ADRG, IDSELI;
output PSADO31, PSADO30, PSADO29, PSADO28, PSADO27, PSADO26, PSADO25, PSADO24, 
    PSADO23, PSADO22, PSADO21, PSADO20, PSADO19, PSADO18, PSADO17, PSADO16, 
    PSADO15, PSADO14, PSADO13, PSADO12, PSADO11, PSADO10, PSADO9, PSADO8, 
    PSADO7, PSADO6, PSADO5, PSADO4, PSADO3, PSADO2, PSADO1, PSADO0, UHIT, 
    ULRDY, CFGW, REGW, REGR, REGADS, RDYACK, LCMD0, ADS, PA7I, PA6I, PA5I, 
    PA4I, PA3I, PA2I;
    wire XADR_30, XADR_17, SPAREO6, LIDSEL, XADR_22, XADR_25, SPAREO0_, 
        SPAREO8, LCMD3, XADR_19, SPAREO1, XADR_10, XADR_18, SPAREO9, XADR_24, 
        XADR_11, SPAREO0, LCMD2, SPAREO7, XADR_31, XADR_16, XADR_23, HitIOL, 
        LAD8, XADR_14, SPAREO5, XADR_28, LAD1, IORCYCA, XADR_21, XADR_26, 
        XADR_8, SPAREO2, XADR_13, XADR_9, HitIOH, XADR_27, XADR_12, SPAREO3, 
        SPAREO1_, LCMD1, XADR_29, IORCYC, SPAREO4, LAD10, LAD9, XADR_15, 
        XADR_20, IOWCYC, LAD0, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
        n1439, n1440, net36, net39, net43, net46, net63, net74, n1441, n1442, 
        n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
        n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
        n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
        n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
        n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
        n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
        n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
        n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520;
    zaoi211b SPARE732 ( .A(SPAREO0), .B(IOWCYC), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE735 ( .A(SPAREO1), .B(HitIOL), .C(SPAREO9), .Y(SPAREO3) );
    zoai21b SPARE734 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE733 ( .A(SPAREO4), .B(HitIOH), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zan2b DNTADS ( .A(UADS), .B(EN_EHCI), .Y(ADS) );
    zdffrb SPARE731 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE738 ( .A(SPAREO5), .Y(SPAREO6) );
    znr3b SPARE736 ( .A(SPAREO2), .B(IORCYCA), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE737 ( .A(SPAREO4), .Y(SPAREO5) );
    zdffrb SPARE730 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE739 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zbfb drv1 ( .A(IORCYCA), .Y(IORCYC) );
    zymx24hb U96 ( .A1(CFGD3), .A2(CFGD2), .A3(CFGD1), .A4(CFGD0), .B1(REGD3), 
        .B2(REGD2), .B3(REGD1), .B4(REGD0), .S(IORCYC), .Y1(PSADO3), .Y2(
        PSADO2), .Y3(PSADO1), .Y4(PSADO0) );
    zymx24hb U97 ( .A1(CFGD7), .A2(CFGD6), .A3(CFGD5), .A4(CFGD4), .B1(REGD7), 
        .B2(REGD6), .B3(REGD5), .B4(REGD4), .S(IORCYC), .Y1(PSADO7), .Y2(
        PSADO6), .Y3(PSADO5), .Y4(PSADO4) );
    zymx24hb U98 ( .A1(CFGD11), .A2(CFGD10), .A3(CFGD9), .A4(CFGD8), .B1(
        REGD11), .B2(REGD10), .B3(REGD9), .B4(REGD8), .S(IORCYC), .Y1(PSADO11), 
        .Y2(PSADO10), .Y3(PSADO9), .Y4(PSADO8) );
    zymx24hb U99 ( .A1(CFGD15), .A2(CFGD14), .A3(CFGD13), .A4(CFGD12), .B1(
        REGD15), .B2(REGD14), .B3(REGD13), .B4(REGD12), .S(IORCYC), .Y1(
        PSADO15), .Y2(PSADO14), .Y3(PSADO13), .Y4(PSADO12) );
    zymx24hb U100 ( .A1(CFGD19), .A2(CFGD18), .A3(CFGD17), .A4(CFGD16), .B1(
        REGD19), .B2(REGD18), .B3(REGD17), .B4(REGD16), .S(IORCYC), .Y1(
        PSADO19), .Y2(PSADO18), .Y3(PSADO17), .Y4(PSADO16) );
    zymx24hb U101 ( .A1(CFGD23), .A2(CFGD22), .A3(CFGD21), .A4(CFGD20), .B1(
        REGD23), .B2(REGD22), .B3(REGD21), .B4(REGD20), .S(IORCYC), .Y1(
        PSADO23), .Y2(PSADO22), .Y3(PSADO21), .Y4(PSADO20) );
    zymx24hb U102 ( .A1(CFGD27), .A2(CFGD26), .A3(CFGD25), .A4(CFGD24), .B1(
        REGD27), .B2(REGD26), .B3(REGD25), .B4(REGD24), .S(IORCYC), .Y1(
        PSADO27), .Y2(PSADO26), .Y3(PSADO25), .Y4(PSADO24) );
    zymx24hb U103 ( .A1(CFGD31), .A2(CFGD30), .A3(CFGD29), .A4(CFGD28), .B1(
        REGD31), .B2(REGD30), .B3(REGD29), .B4(REGD28), .S(IORCYC), .Y1(
        PSADO31), .Y2(PSADO30), .Y3(PSADO29), .Y4(PSADO28) );
    zxn2b U104 ( .A(XADR_20), .B(IOBA20), .Y(n1517) );
    zxn2b U105 ( .A(XADR_27), .B(IOBA27), .Y(n1516) );
    zxn2b U106 ( .A(XADR_22), .B(IOBA22), .Y(n1515) );
    zxn2b U107 ( .A(XADR_21), .B(IOBA21), .Y(n1514) );
    zxn2b U108 ( .A(XADR_19), .B(IOBA19), .Y(n1513) );
    zxn2b U109 ( .A(XADR_16), .B(IOBA16), .Y(n1512) );
    zxn2b U110 ( .A(XADR_28), .B(IOBA28), .Y(n1511) );
    zxn2b U111 ( .A(XADR_18), .B(IOBA18), .Y(n1510) );
    zxo2b U112 ( .A(XADR_26), .B(IOBA26), .Y(n1504) );
    zxo2b U113 ( .A(XADR_31), .B(IOBA31), .Y(n1503) );
    zxo2b U114 ( .A(XADR_29), .B(IOBA29), .Y(n1506) );
    zxo2b U115 ( .A(XADR_23), .B(IOBA23), .Y(n1505) );
    zxn2b U116 ( .A(XADR_12), .B(IOBA12), .Y(n1494) );
    zxn2b U117 ( .A(XADR_15), .B(IOBA15), .Y(n1493) );
    zxn2b U118 ( .A(XADR_13), .B(IOBA13), .Y(n1492) );
    zxn2b U119 ( .A(XADR_8), .B(IOBA8), .Y(n1491) );
    zxn2b U120 ( .A(IOBA14), .B(XADR_14), .Y(n1490) );
    zxn2b U121 ( .A(IOBA9), .B(XADR_9), .Y(n1489) );
    zxn2b U122 ( .A(IOBA11), .B(XADR_11), .Y(n1488) );
    zxn2b U123 ( .A(IOBA10), .B(XADR_10), .Y(n1487) );
    znd5b U124 ( .A(LCMD3), .B(LIDSEL), .C(n1507), .D(n1508), .E(n1509), .Y(
        n1502) );
    zxn2b U125 ( .A(LAD9), .B(FUNCSEL[1]), .Y(n1507) );
    zxn2b U126 ( .A(LAD10), .B(FUNCSEL[2]), .Y(n1508) );
    zxn2b U127 ( .A(LAD8), .B(FUNCSEL[0]), .Y(n1509) );
    zxo2b U128 ( .A(XADR_25), .B(IOBA25), .Y(n1481) );
    zxo2b U129 ( .A(XADR_17), .B(IOBA17), .Y(n1482) );
    zxo2b U130 ( .A(XADR_24), .B(IOBA24), .Y(n1483) );
    zxo2b U131 ( .A(XADR_30), .B(IOBA30), .Y(n1484) );
    znd8b U132 ( .A(n1510), .B(n1511), .C(n1512), .D(n1513), .E(n1514), .F(
        n1515), .G(n1516), .H(n1517), .Y(n1486) );
    zivb U133 ( .A(HitIOL), .Y(n1519) );
    znd8b U134 ( .A(n1487), .B(n1488), .C(n1489), .D(n1490), .E(n1491), .F(
        n1492), .G(n1493), .H(n1494), .Y(HitIOL) );
    zmux21hb U135 ( .A(XADR_16), .B(AD16I), .S(n1438), .Y(n1441) );
    zmux21lb U136 ( .A(net36), .B(n1436), .S(n1439), .Y(n1442) );
    zmux21hb U137 ( .A(LCMD0), .B(CBE0I_), .S(n1438), .Y(n1443) );
    zmux21hb U138 ( .A(XADR_24), .B(AD24I), .S(n1438), .Y(n1444) );
    zmux21lb U139 ( .A(net39), .B(n1437), .S(n1439), .Y(n1445) );
    zmux21hb U140 ( .A(PA7I), .B(AD7I), .S(n1438), .Y(n1446) );
    zmux21hb U141 ( .A(XADR_19), .B(AD19I), .S(n1438), .Y(n1447) );
    zmux21hb U142 ( .A(XADR_22), .B(AD22I), .S(ADRG), .Y(n1448) );
    zmux21lb U143 ( .A(net43), .B(n1435), .S(n1438), .Y(n1449) );
    zmux21hb U144 ( .A(XADR_17), .B(AD17I), .S(n1439), .Y(n1450) );
    zmux21hb U145 ( .A(XADR_25), .B(AD25I), .S(ADRG), .Y(n1451) );
    zmux21lb U146 ( .A(net46), .B(n1436), .S(n1439), .Y(n1452) );
    zivb U147 ( .A(AD8I), .Y(n1436) );
    zmux21hb U148 ( .A(XADR_11), .B(AD11I), .S(ADRG), .Y(n1453) );
    zmux21hb U149 ( .A(XADR_23), .B(AD23I), .S(ADRG), .Y(n1454) );
    zmux21hb U150 ( .A(PA6I), .B(AD6I), .S(n1439), .Y(n1455) );
    zmux21hb U151 ( .A(XADR_18), .B(AD18I), .S(n1439), .Y(n1456) );
    zmux21hb U152 ( .A(LAD0), .B(AD0I), .S(n1439), .Y(n1457) );
    zmux21hb U153 ( .A(LCMD2), .B(CBE2I_), .S(n1439), .Y(n1458) );
    zmux21hb U154 ( .A(PA2I), .B(AD2I), .S(n1439), .Y(n1459) );
    zmux21hb U155 ( .A(XADR_27), .B(AD27I), .S(n1439), .Y(n1460) );
    zmux21hb U156 ( .A(LIDSEL), .B(IDSELI), .S(n1439), .Y(n1461) );
    zmux21hb U157 ( .A(XADR_31), .B(AD31I), .S(n1438), .Y(n1462) );
    zmux21hb U158 ( .A(LAD1), .B(AD1I), .S(n1439), .Y(n1463) );
    zmux21hb U159 ( .A(XADR_15), .B(AD15I), .S(n1438), .Y(n1464) );
    zmux21hb U160 ( .A(XADR_21), .B(AD21I), .S(n1439), .Y(n1465) );
    zmux21hb U161 ( .A(PA4I), .B(AD4I), .S(ADRG), .Y(n1466) );
    zmux21hb U162 ( .A(XADR_28), .B(AD28I), .S(n1439), .Y(n1467) );
    zmux21hb U163 ( .A(XADR_13), .B(AD13I), .S(ADRG), .Y(n1468) );
    zmux21lb U164 ( .A(net63), .B(n1437), .S(n1438), .Y(n1469) );
    zivb U165 ( .A(AD10I), .Y(n1437) );
    zmux21hb U166 ( .A(LCMD3), .B(CBE3I_), .S(n1439), .Y(n1470) );
    zmux21hb U167 ( .A(XADR_26), .B(AD26I), .S(ADRG), .Y(n1471) );
    zmux21hb U168 ( .A(PA3I), .B(AD3I), .S(ADRG), .Y(n1472) );
    zmux21hb U169 ( .A(XADR_14), .B(AD14I), .S(n1439), .Y(n1473) );
    zmux21hb U170 ( .A(XADR_30), .B(AD30I), .S(n1438), .Y(n1474) );
    zmux21hb U171 ( .A(PA5I), .B(AD5I), .S(n1438), .Y(n1475) );
    zmux21hb U172 ( .A(XADR_20), .B(AD20I), .S(n1438), .Y(n1476) );
    zmux21hb U173 ( .A(XADR_12), .B(AD12I), .S(n1438), .Y(n1477) );
    zmux21hb U174 ( .A(XADR_29), .B(AD29I), .S(n1438), .Y(n1478) );
    zmux21hb U175 ( .A(LCMD1), .B(CBE1I_), .S(n1438), .Y(n1479) );
    zmux21lb U176 ( .A(net74), .B(n1435), .S(n1438), .Y(n1480) );
    zivb U177 ( .A(AD9I), .Y(n1435) );
    znr2b U178 ( .A(IRDYI_), .B(TRDYI_), .Y(RDYACK) );
    zor2b U179 ( .A(REGR), .B(REGW), .Y(REGADS) );
    zivb U180 ( .A(IORCYC), .Y(n1501) );
    zivb U181 ( .A(n1500), .Y(IOWCYC) );
    zan3b U182 ( .A(ADS), .B(LCMD0), .C(n1495), .Y(CFGW) );
    zan2b U183 ( .A(ADS), .B(UHIT), .Y(ULRDY) );
    zivb U184 ( .A(ADS), .Y(n1499) );
    znd4b U185 ( .A(IOSPACE), .B(EN_EHCI), .C(n1520), .D(n1518), .Y(n1497) );
    zivb U186 ( .A(HitIOH), .Y(n1520) );
    zivb U187 ( .A(EN_EHCI), .Y(n1496) );
    zivb U188 ( .A(n1498), .Y(n1495) );
    zoa211b U189 ( .A(LCMD1), .B(LCMD3), .C(LCMD2), .D(n1434), .Y(IORCYCA) );
    znr2b U190 ( .A(n1499), .B(n1500), .Y(REGW) );
    znr2b U191 ( .A(n1499), .B(n1501), .Y(REGR) );
    zaoi21b U192 ( .A(n1497), .B(n1498), .C(PMSTR), .Y(UHIT) );
    zivb U193 ( .A(ADRG), .Y(n1440) );
    zivc U194 ( .A(n1440), .Y(n1439) );
    zivc U195 ( .A(n1440), .Y(n1438) );
    zdffb PA16I_reg ( .CK(PCICLK), .D(n1441), .Q(XADR_16) );
    zdffb PA8I_reg ( .CK(PCICLK), .D(n1442), .Q(XADR_8), .QN(net36) );
    zdffb LCMD0_reg ( .CK(PCICLK), .D(n1443), .Q(LCMD0), .QN(n1434) );
    zdffb PA24I_reg ( .CK(PCICLK), .D(n1444), .Q(XADR_24) );
    zdffb PA10I_reg ( .CK(PCICLK), .D(n1445), .Q(XADR_10), .QN(net39) );
    zdffb PA7I_reg ( .CK(PCICLK), .D(n1446), .Q(PA7I) );
    zdffb PA19I_reg ( .CK(PCICLK), .D(n1447), .Q(XADR_19) );
    zdffb PA22I_reg ( .CK(PCICLK), .D(n1448), .Q(XADR_22) );
    zdffb PA9I_reg ( .CK(PCICLK), .D(n1449), .Q(XADR_9), .QN(net43) );
    zdffb PA17I_reg ( .CK(PCICLK), .D(n1450), .Q(XADR_17) );
    zdffb PA25I_reg ( .CK(PCICLK), .D(n1451), .Q(XADR_25) );
    zdffb LAD8_reg ( .CK(PCICLK), .D(n1452), .Q(LAD8), .QN(net46) );
    zdffb PA11I_reg ( .CK(PCICLK), .D(n1453), .Q(XADR_11) );
    zdffb PA23I_reg ( .CK(PCICLK), .D(n1454), .Q(XADR_23) );
    zdffb PA6I_reg ( .CK(PCICLK), .D(n1455), .Q(PA6I) );
    zdffb PA18I_reg ( .CK(PCICLK), .D(n1456), .Q(XADR_18) );
    zdffb LAD0_reg ( .CK(PCICLK), .D(n1457), .Q(LAD0) );
    zdffb LCMD2_reg ( .CK(PCICLK), .D(n1458), .Q(LCMD2), .QN(n1433) );
    zdffb PA2I_reg ( .CK(PCICLK), .D(n1459), .Q(PA2I) );
    zdffb PA27I_reg ( .CK(PCICLK), .D(n1460), .Q(XADR_27) );
    zdffb LIDSEL_reg ( .CK(PCICLK), .D(n1461), .Q(LIDSEL) );
    zdffb PA31I_reg ( .CK(PCICLK), .D(n1462), .Q(XADR_31) );
    zdffb LAD1_reg ( .CK(PCICLK), .D(n1463), .Q(LAD1) );
    zdffb PA15I_reg ( .CK(PCICLK), .D(n1464), .Q(XADR_15) );
    zdffb PA21I_reg ( .CK(PCICLK), .D(n1465), .Q(XADR_21) );
    zdffb PA4I_reg ( .CK(PCICLK), .D(n1466), .Q(PA4I) );
    zdffb PA28I_reg ( .CK(PCICLK), .D(n1467), .Q(XADR_28) );
    zdffb PA13I_reg ( .CK(PCICLK), .D(n1468), .Q(XADR_13) );
    zdffb LAD10_reg ( .CK(PCICLK), .D(n1469), .Q(LAD10), .QN(net63) );
    zdffb LCMD3_reg ( .CK(PCICLK), .D(n1470), .Q(LCMD3) );
    zdffb PA26I_reg ( .CK(PCICLK), .D(n1471), .Q(XADR_26) );
    zdffb PA3I_reg ( .CK(PCICLK), .D(n1472), .Q(PA3I) );
    zdffb PA14I_reg ( .CK(PCICLK), .D(n1473), .Q(XADR_14) );
    zdffb PA30I_reg ( .CK(PCICLK), .D(n1474), .Q(XADR_30) );
    zdffb PA5I_reg ( .CK(PCICLK), .D(n1475), .Q(PA5I) );
    zdffb PA20I_reg ( .CK(PCICLK), .D(n1476), .Q(XADR_20) );
    zdffb PA12I_reg ( .CK(PCICLK), .D(n1477), .Q(XADR_12) );
    zdffb PA29I_reg ( .CK(PCICLK), .D(n1478), .Q(XADR_29) );
    zdffb LCMD1_reg ( .CK(PCICLK), .D(n1479), .Q(LCMD1), .QN(n1432) );
    zdffb LAD9_reg ( .CK(PCICLK), .D(n1480), .Q(LAD9), .QN(net74) );
    zor6b U196 ( .A(n1481), .B(n1482), .C(n1483), .D(n1484), .E(n1485), .F(
        n1486), .Y(HitIOH) );
    zor3b U197 ( .A(n1432), .B(n1433), .C(n1434), .Y(n1500) );
    zor6b U198 ( .A(LAD1), .B(LAD0), .C(LCMD2), .D(n1432), .E(n1496), .F(n1502
        ), .Y(n1498) );
    zor4b U199 ( .A(n1505), .B(n1506), .C(n1503), .D(n1504), .Y(n1485) );
    zoa21d U200 ( .A(IOWCYC), .B(IORCYC), .C(n1519), .Y(n1518) );
endmodule


module HS_OPREG ( REGD31, REGD30, REGD29, REGD28, REGD27, REGD26, REGD25, 
    REGD24, REGD23, REGD22, REGD21, REGD20, REGD19, REGD18, REGD17, REGD16, 
    REGD15, REGD14, REGD13, REGD12, REGD11, REGD10, REGD9, REGD8, REGD7, REGD6, 
    REGD5, REGD4, REGD3, REGD2, REGD1, REGD0, REGDOUT2, LIGHTRST, INTDOORBELL, 
    ASYNC_EN, PERIOD_EN, HCRESET, RUN, INTTHRESHOLD, FRLSTSIZE, MABORTS, 
    TABORTR, RUN_C, INTASYNC_EN, HSERR_EN, ROLLOVER_EN, PORTCHG_EN, ERRINT_EN, 
    USBINT_EN, FLBASE, ASYNCLISTADDR, WR_FRNUM, WR_ASYNCADDR, USBINT, ERRINT, 
    INTASYNC, ASYNCINT, UINTOE_, HCHALT, CMDRST_, HSERR_S, DBGIRQ, UIRQACT, 
    USBLEGCTLSTS, USBLEGSUP, USMIO, ASYNC_ACT, PERIOD_ACT, RECLAMATION, 
    MAC_EOT, EHCI_IDLE, INTASYNC_S, ROLLOVER_S, PORTCHG_S, ERRINT_S, USBINT_S, 
    PWR_STATE_D0, PORTSC1, PORTSC2, PORTSC3, PORTSC4, PORTSC5, PORTSC6, 
    PORTSC7, PORTSC8, CFG_CS, PSC_CBE2_A, PSC_CBE1_A, PSC_CBE0_A, PSC_CBE2_B, 
    PSC_CBE1_B, PSC_CBE0_B, PSC_CBE2_C, PSC_CBE1_C, PSC_CBE0_C, PSC_CBE2_D, 
    PSC_CBE1_D, PSC_CBE0_D, PSC_CBE2_E, PSC_CBE1_E, PSC_CBE0_E, PSC_CBE2_F, 
    PSC_CBE1_F, PSC_CBE0_F, PSC_CBE2_G, PSC_CBE1_G, PSC_CBE0_G, PSC_CBE2_H, 
    PSC_CBE1_H, PSC_CBE0_H, AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, 
    AD24I, AD23I, AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, 
    AD14I, AD13I, AD12I, AD11I, AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, 
    AD3I, AD2I, AD1I, AD0I, CBE3I_, CBE2I_, CBE1I_, CBE0I_, REGW, PA7I, PA6I, 
    PA5I, PA4I, PA3I, PA2I, FRNUM, FRNUM_PCLK_LATCH_66, ConfigFlag, 
    TEST_FORCE_ENABLE, PCI_R6AG, PCI_R6BG, PCI_R6CG, PCI_R6DG, PCI_R6FG, 
    PCI_RBAR, PCI_RPCMD, INTR_DIS, SUBIDWE, PCICLK, PCICLK_FREE, HRST_, 
    ATPG_ENI, ENUSB1, ENUSB2, ENUSB3, ENUSB4, DIS_SOF_RUN, UTM_RUN, 
    EN_DBG_PORT, DBGPORT_R00G, DBGPORT_R01G, DBGPORT_R02G, DBGPORT_R03G, 
    DBGPORT_R04G, DBGPORT_R05G, DBGPORT_R08G, DBGPORT_R09G, DBGPORT_R0AG, 
    DBGPORT_R0BG, DBGPORT_R0CG, DBGPORT_R0DG, DBGPORT_R0EG, DBGPORT_R0FG, 
    DBGPORT_R10G, DBGPORT_R11G, DBGPORT_SC, DBGPORT_PID, DBGPORT_ADDR, 
    DBGPORT_BUF1, DBGPORT_BUF2 );
output [31:0] REGDOUT2;
output [1:0] FRLSTSIZE;
input  [31:0] PORTSC7;
input  [31:0] PORTSC6;
input  [13:0] FRNUM;
input  [31:0] PORTSC8;
input  [31:0] DBGPORT_BUF2;
output [7:0] INTTHRESHOLD;
input  [31:0] ASYNCLISTADDR;
output [31:0] USBLEGSUP;
input  [31:0] PORTSC1;
input  [31:0] PORTSC3;
output [31:12] FLBASE;
input  [31:0] PORTSC4;
input  [31:0] DBGPORT_SC;
input  [31:0] DBGPORT_PID;
output [31:0] USBLEGCTLSTS;
input  [31:0] PORTSC2;
input  [31:0] PORTSC5;
input  [31:0] DBGPORT_ADDR;
input  [31:0] DBGPORT_BUF1;
input  MABORTS, TABORTR, RUN_C, ASYNCINT, HSERR_S, DBGIRQ, ASYNC_ACT, 
    PERIOD_ACT, RECLAMATION, MAC_EOT, EHCI_IDLE, INTASYNC_S, ROLLOVER_S, 
    PORTCHG_S, ERRINT_S, USBINT_S, PWR_STATE_D0, AD31I, AD30I, AD29I, AD28I, 
    AD27I, AD26I, AD25I, AD24I, AD23I, AD22I, AD21I, AD20I, AD19I, AD18I, 
    AD17I, AD16I, AD15I, AD14I, AD13I, AD12I, AD11I, AD10I, AD9I, AD8I, AD7I, 
    AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I, CBE3I_, CBE2I_, CBE1I_, CBE0I_, 
    REGW, PA7I, PA6I, PA5I, PA4I, PA3I, PA2I, FRNUM_PCLK_LATCH_66, ConfigFlag, 
    TEST_FORCE_ENABLE, PCI_R6AG, PCI_R6BG, PCI_R6CG, PCI_R6DG, PCI_R6FG, 
    PCI_RBAR, PCI_RPCMD, INTR_DIS, SUBIDWE, PCICLK, PCICLK_FREE, HRST_, 
    ATPG_ENI, ENUSB1, ENUSB2, ENUSB3, ENUSB4, DIS_SOF_RUN, EN_DBG_PORT;
output REGD31, REGD30, REGD29, REGD28, REGD27, REGD26, REGD25, REGD24, REGD23, 
    REGD22, REGD21, REGD20, REGD19, REGD18, REGD17, REGD16, REGD15, REGD14, 
    REGD13, REGD12, REGD11, REGD10, REGD9, REGD8, REGD7, REGD6, REGD5, REGD4, 
    REGD3, REGD2, REGD1, REGD0, LIGHTRST, INTDOORBELL, ASYNC_EN, PERIOD_EN, 
    HCRESET, RUN, INTASYNC_EN, HSERR_EN, ROLLOVER_EN, PORTCHG_EN, ERRINT_EN, 
    USBINT_EN, WR_FRNUM, WR_ASYNCADDR, USBINT, ERRINT, INTASYNC, UINTOE_, 
    HCHALT, CMDRST_, UIRQACT, USMIO, CFG_CS, PSC_CBE2_A, PSC_CBE1_A, 
    PSC_CBE0_A, PSC_CBE2_B, PSC_CBE1_B, PSC_CBE0_B, PSC_CBE2_C, PSC_CBE1_C, 
    PSC_CBE0_C, PSC_CBE2_D, PSC_CBE1_D, PSC_CBE0_D, PSC_CBE2_E, PSC_CBE1_E, 
    PSC_CBE0_E, PSC_CBE2_F, PSC_CBE1_F, PSC_CBE0_F, PSC_CBE2_G, PSC_CBE1_G, 
    PSC_CBE0_G, PSC_CBE2_H, PSC_CBE1_H, PSC_CBE0_H, UTM_RUN, DBGPORT_R00G, 
    DBGPORT_R01G, DBGPORT_R02G, DBGPORT_R03G, DBGPORT_R04G, DBGPORT_R05G, 
    DBGPORT_R08G, DBGPORT_R09G, DBGPORT_R0AG, DBGPORT_R0BG, DBGPORT_R0CG, 
    DBGPORT_R0DG, DBGPORT_R0EG, DBGPORT_R0FG, DBGPORT_R10G, DBGPORT_R11G;
    wire n_561, HCSPARAMS_9, n_1886, HCRESET1670, SPAREO6, SMIHERR_EN2413, 
        HCIVERSION_3, FRNUM_SYNC_8, RAEG, INTTHRESHOLD1414_1, n_1878, 
        HCSPARAMS_12, n_834, val1944_1, HCIVERSION_10, HCSPARAMS_0, 
        FLBASE2087_19, n_1240, ENUSB_1, FRNUM_SYNC_1, PORTCHG_EN1992, RAAG, 
        FLBASE2087_25, FRNUM_SYNC_13, LIGHTRST_2T, n_1876, HCRESET_2T, RACG, 
        FLBASE2087_22, ERRINT_EN1986, HCCPARAMS_4, FRNUM_SYNC_6, SPAREO0_, 
        OSOWNS2125, n_1888, SPAREO8, n_1613, PERIOD_STS, USMIO_2T, HCSPARAMS_7, 
        SMIONPCMD_EN2320, n_1601, INTTHRESHOLD1414_6, n_2155, HCCPARAMS_13, 
        SPAREO1, n_846, FLBASE2087_30, FLBASE2087_17, USBSTS1, HCSPARAMS_6, 
        n_2161, n_1246, SPAREO9, FRNUM_SYNC_7, HSERR_EN2004, FLBASE2087_23, 
        n_1609, HCCPARAMS_5, BIOSOWNS2162, FLBASE2087_31, n_567, FLBASE2087_16, 
        USBSTS0, USBSMI_EN2389, n_1880, USMIACT_T, SPAREO0, HCIVERSION_5, 
        INTTHRESHOLD1414_7, HCSPARAMS_14, SMIPORTCHG_EN2401, n_832, 
        HCSPARAMS_13, n_1607, RA8G, PERIOD_EN1619, HCIVERSION_2, FRNUM_SYNC_9, 
        INTTHRESHOLD1414_0, n_2153, n_840, n_1248, SPAREO7, INTASYNC_EN2010, 
        SMIOWN_EN2314, ROLLOVER_EN1998, HCSPARAMS_8, FLBASE2087_24, 
        FRNUM_SYNC_12, UTM_RUN_T, FRNUM_SYNC_0, ASYNC_STS, ENUSB_0, n_1615, 
        HCIVERSION_11, HCSPARAMS_1, n_569, FLBASE2087_18, USBSTS5, 
        FLBASE2087_13, n_842, SPAREO5, n_15, n_2151, INTTHRESHOLD1414_2, 
        HCIVERSION_0, n_1605, HCCPARAMS_9, HCSPARAMS_11, RA9G, HCSPARAMS_3, 
        HCIVERSION_13, SMIONBAR_NXT, n3526, ENUSB_2, RUN1760, USBINT_EN1980, 
        FRNUM_SYNC_2, HCIVERSION_9, HCCPARAMS_0, n_557, FLBASE2087_26, USMIACT, 
        FRNUM_SYNC_10, n_1236, HCCPARAMS_7, INTDOORBELL1489, USMIO_T2541, 
        FLBASE2087_21, n_1890, FRNUM_SYNC_5, n_1244, LIGHTRST1452, n_2163, 
        HCSPARAMS_4, HCIVERSION_14, n_12, n_559, FLBASE2087_28, n_1238, 
        FRLSTSIZE1579_1, n_3593, INTTHRESHOLD1414_5, HCIVERSION_7, n_1882, 
        SPAREO2, HCCPARAMS_10, SMIUSBERR_EN2395, FLBASE2087_14, n_565, USBSTS2, 
        HCRESET_T, HCSPARAMS_5, HCIVERSION_15, n_1611, val1876_1, RAFG, 
        USMIO_T, SMIFROVER_EN2407, FRNUM_SYNC_4, HCCPARAMS_6, ASYNC_EN1625, 
        n_838, RABG, FLBASE2087_20, FLBASE2087_15, USBSTS3, REGX0, SPAREO3, 
        n_844, SMIONPCMD_NXT, HCCPARAMS_11, SPAREO1_, n_2157, 
        INTTHRESHOLD1414_4, n_13, HCIVERSION_6, n_1603, FLBASE2087_29, 
        LIGHTRST_T, USMIO_3T, FRLSTSIZE1579_0, HCCPARAMS_8, n_14, n_836, 
        HCSPARAMS_10, n_1250, INTTHRESHOLD1414_3, HCIVERSION_1, 
        SMIOSOWNCHG_NXT, n_1884, SPAREO4, SMIONBAR_EN2326, USBSTS4, 
        FLBASE2087_12, n_563, FLBASE2087_27, FRNUM_SYNC_11, n_571, 
        SMIASYNC_EN2419, n_2159, FRNUM_SYNC_3, HCIVERSION_8, ENUSB_3, n_2165, 
        RADG, n_1242, HCSPARAMS_2, HCIVERSION_12, n2977, n2978, n2979, n2980, 
        n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, 
        n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
        n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, 
        n3011, n3012, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
        n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
        n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
        n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
        n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
        n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
        n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
        n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
        n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
        n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
        n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
        n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
        n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
        n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
        n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
        n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, 
        n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
        n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
        n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, 
        n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, 
        n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, 
        n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
        n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, 
        n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, 
        n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, 
        n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, 
        n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, 
        n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, 
        n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, 
        n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, 
        n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, 
        n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, 
        n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, 
        n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, 
        n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, 
        n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, 
        n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, 
        n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, 
        n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, 
        n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, 
        n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, 
        n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, 
        n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, 
        n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, 
        n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, 
        n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, 
        n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, 
        n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, 
        n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, 
        n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, 
        n3514, n3517, n3518, n3519, n3520, n3521, n3522, n3524, n3525;
    assign USBLEGCTLSTS[28] = 1'b0;
    assign USBLEGCTLSTS[27] = 1'b0;
    assign USBLEGCTLSTS[26] = 1'b0;
    assign USBLEGCTLSTS[25] = 1'b0;
    assign USBLEGCTLSTS[24] = 1'b0;
    assign USBLEGCTLSTS[23] = 1'b0;
    assign USBLEGCTLSTS[22] = 1'b0;
    assign USBLEGCTLSTS[12] = 1'b0;
    assign USBLEGCTLSTS[11] = 1'b0;
    assign USBLEGCTLSTS[10] = 1'b0;
    assign USBLEGCTLSTS[9] = 1'b0;
    assign USBLEGCTLSTS[8] = 1'b0;
    assign USBLEGCTLSTS[7] = 1'b0;
    assign USBLEGCTLSTS[6] = 1'b0;
    assign USBLEGSUP[31] = 1'b0;
    assign USBLEGSUP[30] = 1'b0;
    assign USBLEGSUP[29] = 1'b0;
    assign USBLEGSUP[28] = 1'b0;
    assign USBLEGSUP[27] = 1'b0;
    assign USBLEGSUP[26] = 1'b0;
    assign USBLEGSUP[25] = 1'b0;
    assign USBLEGSUP[23] = 1'b0;
    assign USBLEGSUP[22] = 1'b0;
    assign USBLEGSUP[21] = 1'b0;
    assign USBLEGSUP[20] = 1'b0;
    assign USBLEGSUP[19] = 1'b0;
    assign USBLEGSUP[18] = 1'b0;
    assign USBLEGSUP[17] = 1'b0;
    assign USBLEGSUP[15] = 1'b0;
    assign USBLEGSUP[14] = 1'b0;
    assign USBLEGSUP[13] = 1'b0;
    assign USBLEGSUP[12] = 1'b0;
    assign USBLEGSUP[11] = 1'b0;
    assign USBLEGSUP[10] = 1'b0;
    assign USBLEGSUP[9] = 1'b0;
    assign USBLEGSUP[8] = 1'b0;
    assign USBLEGSUP[7] = 1'b0;
    assign USBLEGSUP[6] = 1'b0;
    assign USBLEGSUP[5] = 1'b0;
    assign USBLEGSUP[4] = 1'b0;
    assign USBLEGSUP[3] = 1'b0;
    assign USBLEGSUP[2] = 1'b0;
    assign USBLEGSUP[1] = 1'b0;
    assign USBLEGSUP[0] = 1'b1;
    zivb SPARE747 ( .A(SPAREO4), .Y(SPAREO5) );
    znd3b SPARE749 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE740 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE748 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE741 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    znr3b SPARE746 ( .A(SPAREO2), .B(REGX0), .C(SPAREO0_), .Y(SPAREO4) );
    zoai21b SPARE744 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE743 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zaoi211b SPARE742 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE745 ( .A(SPAREO1), .B(SMIONBAR_NXT), .C(SPAREO9), .Y(SPAREO3)
         );
    zao33b U718 ( .A(USBLEGCTLSTS[15]), .B(n3347), .C(SMIONBAR_NXT), .D(
        USBLEGCTLSTS[5]), .E(n3357), .F(INTASYNC_S), .Y(n3033) );
    zao33b U719 ( .A(USBLEGCTLSTS[1]), .B(n3355), .C(USBSTS1), .D(USBLEGCTLSTS
        [3]), .E(n3353), .F(USBSTS3), .Y(n3031) );
    zao33b U720 ( .A(USBLEGCTLSTS[4]), .B(n3351), .C(USBSTS4), .D(USBLEGCTLSTS
        [2]), .E(n3349), .F(USBSTS2), .Y(n3030) );
    zivb U721 ( .A(ENUSB1), .Y(n3255) );
    zivb U722 ( .A(ENUSB3), .Y(n3256) );
    zxo2b U723 ( .A(ENUSB_3), .B(ENUSB4), .Y(n3324) );
    zxo2b U724 ( .A(ENUSB_2), .B(ENUSB3), .Y(n3325) );
    zxo2b U725 ( .A(ENUSB_0), .B(ENUSB1), .Y(n3326) );
    zxo2b U726 ( .A(ENUSB_1), .B(ENUSB2), .Y(n3327) );
    zor2b U727 ( .A(n3332), .B(n3338), .Y(n3259) );
    zor2b U728 ( .A(PA7I), .B(n3335), .Y(n3336) );
    zao22b U729 ( .A(USBINT_EN), .B(USBINT), .C(ERRINT_EN), .D(ERRINT), .Y(
        n3065) );
    zor2b U730 ( .A(n3294), .B(n3319), .Y(n3337) );
    zao32b U731 ( .A(ConfigFlag), .B(REGX0), .C(n3053), .D(DBGPORT_BUF1[0]), 
        .E(n3513), .Y(n3500) );
    zoai2x4b U732 ( .A(n_12), .B(n3391), .C(n3355), .D(n3394), .E(n3364), .F(
        n3393), .G(n3297), .H(n3312), .Y(n3497) );
    zoai2x4b U733 ( .A(n3349), .B(n3394), .C(n3361), .D(n3393), .E(n3297), .F(
        n3313), .G(n3321), .H(n3333), .Y(n3487) );
    zoai2x4b U734 ( .A(n3353), .B(n3394), .C(n3362), .D(n3393), .E(n3297), .F(
        n3314), .G(n3321), .H(n3334), .Y(n3471) );
    zao22b U735 ( .A(HCCPARAMS_5), .B(n3450), .C(n3458), .D(INTASYNC_EN), .Y(
        n3455) );
    zor2b U736 ( .A(n3295), .B(n3338), .Y(n3393) );
    zoai2x4b U737 ( .A(n3394), .B(n3424), .C(n3321), .D(n3330), .E(n3396), .F(
        n3423), .G(n3297), .H(n3303), .Y(n3495) );
    zao2x4b U738 ( .A(HCSPARAMS_13), .B(n3451), .C(FLBASE[13]), .D(n3465), .E(
        HCCPARAMS_13), .F(n3450), .G(RECLAMATION), .H(n3459), .Y(n3491) );
    zor2b U739 ( .A(n3270), .B(n3295), .Y(n3297) );
    zor2b U740 ( .A(n3320), .B(n3338), .Y(n3394) );
    zor2b U741 ( .A(n3270), .B(n3320), .Y(n3321) );
    zor2b U742 ( .A(n3271), .B(n3338), .Y(n3391) );
    zor2b U743 ( .A(n3369), .B(n3370), .Y(n3371) );
    zor2b U744 ( .A(n3370), .B(n3372), .Y(n3373) );
    zor2b U745 ( .A(n3270), .B(n3271), .Y(n3274) );
    zor2b U746 ( .A(PA5I), .B(n3269), .Y(n3270) );
    zor2b U747 ( .A(PA3I), .B(PA2I), .Y(n3271) );
    zivb U748 ( .A(n3271), .Y(REGX0) );
    zor2b U749 ( .A(PA3I), .B(n3319), .Y(n3320) );
    zivb U750 ( .A(PA2I), .Y(n3319) );
    zor2b U751 ( .A(n3034), .B(INTASYNC_S), .Y(USBSTS5) );
    zor2b U752 ( .A(n3043), .B(ERRINT_S), .Y(USBSTS1) );
    zor2b U753 ( .A(n3036), .B(USBINT_S), .Y(USBSTS0) );
    zmux21hb U754 ( .A(FRNUM_SYNC_13), .B(FRNUM[13]), .S(n_3593), .Y(n3016) );
    zmux21hb U755 ( .A(FRNUM_SYNC_12), .B(FRNUM[12]), .S(n_3593), .Y(n3017) );
    zmux21hb U756 ( .A(FRNUM_SYNC_11), .B(FRNUM[11]), .S(n_3593), .Y(n3018) );
    zmux21hb U757 ( .A(FRNUM_SYNC_10), .B(FRNUM[10]), .S(n_3593), .Y(n3019) );
    zmux21hb U758 ( .A(FRNUM_SYNC_9), .B(FRNUM[9]), .S(n_3593), .Y(n3020) );
    zmux21hb U759 ( .A(FRNUM_SYNC_8), .B(FRNUM[8]), .S(n_3593), .Y(n3021) );
    zmux21hb U760 ( .A(FRNUM_SYNC_7), .B(FRNUM[7]), .S(n_3593), .Y(n3022) );
    zmux21hb U761 ( .A(FRNUM_SYNC_6), .B(FRNUM[6]), .S(n_3593), .Y(n3023) );
    zmux21hb U762 ( .A(FRNUM_SYNC_5), .B(FRNUM[5]), .S(n_3593), .Y(n3024) );
    zmux21hb U763 ( .A(FRNUM_SYNC_4), .B(FRNUM[4]), .S(n_3593), .Y(n3025) );
    zmux21hb U764 ( .A(FRNUM_SYNC_3), .B(FRNUM[3]), .S(n_3593), .Y(n3026) );
    zmux21hb U765 ( .A(FRNUM_SYNC_2), .B(FRNUM[2]), .S(n_3593), .Y(n3027) );
    zmux21hb U766 ( .A(FRNUM_SYNC_1), .B(FRNUM[1]), .S(n_3593), .Y(n3028) );
    zmux21hb U767 ( .A(FRNUM_SYNC_0), .B(FRNUM[0]), .S(n_3593), .Y(n3029) );
    zan2b U768 ( .A(n3054), .B(n3060), .Y(RAFG) );
    zan2b U769 ( .A(n3054), .B(n3055), .Y(RAEG) );
    zan2b U770 ( .A(n3054), .B(n3049), .Y(RADG) );
    zan2b U771 ( .A(n3054), .B(n3051), .Y(RACG) );
    zivb U772 ( .A(n3369), .Y(n3054) );
    zor2b U773 ( .A(n3337), .B(n3368), .Y(n3369) );
    zan2b U774 ( .A(n3052), .B(n3060), .Y(RABG) );
    zan2b U775 ( .A(n3052), .B(n3055), .Y(RAAG) );
    zan2b U776 ( .A(n3052), .B(n3049), .Y(RA9G) );
    zivb U777 ( .A(n3372), .Y(n3052) );
    zor2b U778 ( .A(n3295), .B(n3368), .Y(n3372) );
    zan2b U779 ( .A(n3044), .B(n3066), .Y(RA8G) );
    zivb U780 ( .A(n3264), .Y(n3103) );
    zivb U781 ( .A(n3504), .Y(n3445) );
    zmux21lb U782 ( .A(n3360), .B(n3097), .S(n2977), .Y(HSERR_EN2004) );
    zmux21lb U783 ( .A(n3291), .B(n3436), .S(n2985), .Y(n_561) );
    zmux21lb U784 ( .A(n3280), .B(n3430), .S(n2984), .Y(n_838) );
    zivb U785 ( .A(AD28I), .Y(n3430) );
    zmux21lb U786 ( .A(n3412), .B(n3434), .S(n2978), .Y(INTTHRESHOLD1414_3) );
    zmux21lb U787 ( .A(n3308), .B(n3076), .S(n2986), .Y(n_2151) );
    zmux21lb U788 ( .A(n3440), .B(n3101), .S(n3103), .Y(RUN1760) );
    zcxi4b U789 ( .A(TEST_FORCE_ENABLE), .B(RUN), .C(MABORTS), .D(n3446), .Y(
        n3440) );
    zmux21lb U790 ( .A(n3343), .B(n3304), .S(PCI_R6DG), .Y(SMIOWN_EN2314) );
    zmux21lb U791 ( .A(n3311), .B(n3101), .S(n2987), .Y(n_1890) );
    zor2b U792 ( .A(n3042), .B(PCI_RBAR), .Y(SMIONBAR_NXT) );
    zmux21lb U793 ( .A(n3265), .B(n3097), .S(n3103), .Y(PERIOD_EN1619) );
    zmux21lb U794 ( .A(n3318), .B(n3089), .S(n2987), .Y(n_1876) );
    zmux21lb U795 ( .A(n3303), .B(n3302), .S(n2986), .Y(n_2157) );
    zivb U796 ( .A(AD12I), .Y(n3302) );
    zmux21lb U797 ( .A(n3443), .B(n3093), .S(n3103), .Y(INTDOORBELL1489) );
    zor2b U798 ( .A(INTASYNC_S), .B(n3392), .Y(n3443) );
    zmux21lb U799 ( .A(n3345), .B(n3306), .S(PCI_R6DG), .Y(SMIONPCMD_EN2320)
         );
    zmux21lb U800 ( .A(n3283), .B(n3260), .S(n2984), .Y(n_832) );
    zivb U801 ( .A(AD31I), .Y(n3260) );
    zmux21lb U802 ( .A(n3410), .B(n3435), .S(n2978), .Y(INTTHRESHOLD1414_4) );
    zmux21lb U803 ( .A(n3359), .B(n3101), .S(n2977), .Y(USBINT_EN1980) );
    zmux21lb U804 ( .A(n3288), .B(n3433), .S(n2985), .Y(n_567) );
    zmux21lb U805 ( .A(n3441), .B(n3426), .S(PCI_R6BG), .Y(OSOWNS2125) );
    zmux21lb U806 ( .A(n3305), .B(n3304), .S(n2986), .Y(n_2155) );
    zivb U807 ( .A(AD13I), .Y(n3304) );
    zmux21lb U808 ( .A(n3362), .B(n3109), .S(n2977), .Y(ROLLOVER_EN1998) );
    zmux21lb U809 ( .A(n3317), .B(n3093), .S(n2987), .Y(n_1878) );
    zivb U810 ( .A(AD6I), .Y(n3093) );
    zao21b U811 ( .A(ASYNC_STS), .B(ASYNC_EN), .C(ASYNC_ACT), .Y(val1876_1) );
    zmux21lb U812 ( .A(n3289), .B(n3434), .S(n2985), .Y(n_565) );
    zivb U813 ( .A(AD19I), .Y(n3434) );
    zao21b U814 ( .A(PCI_R6BG), .B(n3037), .C(n3038), .Y(SMIOSOWNCHG_NXT) );
    zxo2b U815 ( .A(USBLEGSUP[24]), .B(AD24I), .Y(n3037) );
    zmux21lb U816 ( .A(n3356), .B(n3261), .S(PCI_R6CG), .Y(SMIUSBERR_EN2395)
         );
    zmux21lb U817 ( .A(n3354), .B(n3109), .S(PCI_R6CG), .Y(SMIFROVER_EN2407)
         );
    zmux21lb U818 ( .A(n3282), .B(n3262), .S(n2984), .Y(n_834) );
    zmux21lb U819 ( .A(n3408), .B(n3436), .S(n2978), .Y(INTTHRESHOLD1414_5) );
    zivb U820 ( .A(AD21I), .Y(n3436) );
    zmux21lb U821 ( .A(n3281), .B(n3257), .S(n2984), .Y(n_836) );
    zivb U822 ( .A(AD29I), .Y(n3257) );
    zmux21lb U823 ( .A(n3414), .B(n3433), .S(n2978), .Y(INTTHRESHOLD1414_2) );
    zivb U824 ( .A(AD18I), .Y(n3433) );
    zor2b U825 ( .A(n3035), .B(PCI_RPCMD), .Y(SMIONPCMD_NXT) );
    zivb U826 ( .A(AD30I), .Y(n3262) );
    zivb U827 ( .A(PCI_R6FG), .Y(n3258) );
    zmux21hb U828 ( .A(USBLEGSUP[16]), .B(AD16I), .S(PCI_R6AG), .Y(
        BIOSOWNS2162) );
    zmux21lb U829 ( .A(n3290), .B(n3435), .S(n2985), .Y(n_563) );
    zivb U830 ( .A(AD20I), .Y(n3435) );
    zmux21lb U831 ( .A(n3363), .B(n3095), .S(n2977), .Y(INTASYNC_EN2010) );
    zmux21lb U832 ( .A(n3312), .B(n3261), .S(n2987), .Y(n_1888) );
    znr2b U833 ( .A(n3518), .B(n3075), .Y(USMIO_T2541) );
    zivb U834 ( .A(USMIACT), .Y(n3075) );
    zmux21lb U835 ( .A(n3307), .B(n3306), .S(n2986), .Y(n_2153) );
    zivb U836 ( .A(AD14I), .Y(n3306) );
    zmux21lb U837 ( .A(n3444), .B(n3261), .S(n3103), .Y(HCRESET1670) );
    zor2b U838 ( .A(HCRESET_2T), .B(n_12), .Y(n3444) );
    zor2b U839 ( .A(n3338), .B(n3366), .Y(n3264) );
    zmux21lb U840 ( .A(n3276), .B(n3426), .S(n2984), .Y(n_846) );
    zivb U841 ( .A(AD24I), .Y(n3426) );
    zmux21lb U842 ( .A(n3267), .B(n3095), .S(n3103), .Y(ASYNC_EN1625) );
    zmux21lb U843 ( .A(n3344), .B(n3101), .S(PCI_R6CG), .Y(USBSMI_EN2389) );
    zivb U844 ( .A(AD0I), .Y(n3101) );
    zmux21lb U845 ( .A(n3292), .B(n3437), .S(n2985), .Y(n_559) );
    zmux21lb U846 ( .A(n3418), .B(n3431), .S(n2978), .Y(INTTHRESHOLD1414_0) );
    zmux21lb U847 ( .A(n3279), .B(n3429), .S(n2984), .Y(n_840) );
    zivb U848 ( .A(AD27I), .Y(n3429) );
    zmux21lb U849 ( .A(n3314), .B(n3109), .S(n2987), .Y(n_1884) );
    zmux21lb U850 ( .A(n3350), .B(n3106), .S(PCI_R6CG), .Y(SMIPORTCHG_EN2401)
         );
    zmux21lb U851 ( .A(n3361), .B(n3106), .S(n2977), .Y(PORTCHG_EN1992) );
    zmux21lb U852 ( .A(n3315), .B(n3097), .S(n2987), .Y(n_1882) );
    zmux21lb U853 ( .A(n3299), .B(n3439), .S(n2986), .Y(n_2163) );
    zmux21lb U854 ( .A(n3301), .B(n3082), .S(n2986), .Y(n_2159) );
    zivb U855 ( .A(AD11I), .Y(n3082) );
    zivb U856 ( .A(ENUSB4), .Y(n3322) );
    zmux21lb U857 ( .A(n3404), .B(n3438), .S(n2978), .Y(INTTHRESHOLD1414_7) );
    zao21b U858 ( .A(PERIOD_STS), .B(PERIOD_EN), .C(PERIOD_ACT), .Y(val1944_1)
         );
    zmux21lb U859 ( .A(n3287), .B(n3432), .S(n2985), .Y(n_569) );
    zmux21lb U860 ( .A(n3348), .B(n3076), .S(PCI_R6DG), .Y(SMIONBAR_EN2326) );
    zmux21lb U861 ( .A(n3346), .B(n3095), .S(PCI_R6CG), .Y(SMIASYNC_EN2419) );
    zmux21lb U862 ( .A(n3298), .B(n3087), .S(n2986), .Y(n_2165) );
    zivb U863 ( .A(AD8I), .Y(n3087) );
    zmux21lb U864 ( .A(n3442), .B(n3089), .S(n3103), .Y(LIGHTRST1452) );
    zor2b U865 ( .A(LIGHTRST_2T), .B(n_14), .Y(n3442) );
    zivb U866 ( .A(AD7I), .Y(n3089) );
    zmux21lb U867 ( .A(n3300), .B(n3084), .S(n2986), .Y(n_2161) );
    zivb U868 ( .A(AD10I), .Y(n3084) );
    zmux21lb U869 ( .A(n3316), .B(n3095), .S(n2987), .Y(n_1880) );
    zivb U870 ( .A(AD5I), .Y(n3095) );
    zmux21lb U871 ( .A(n3286), .B(n3431), .S(n2985), .Y(n_571) );
    zivb U872 ( .A(AD16I), .Y(n3431) );
    zmux21lb U873 ( .A(n3364), .B(n3261), .S(n2977), .Y(ERRINT_EN1986) );
    zivb U874 ( .A(AD1I), .Y(n3261) );
    zmux21lb U875 ( .A(n3352), .B(n3097), .S(PCI_R6CG), .Y(SMIHERR_EN2413) );
    zivb U876 ( .A(n3090), .Y(n3099) );
    zmux21lb U877 ( .A(n3406), .B(n3437), .S(n2978), .Y(INTTHRESHOLD1414_6) );
    zivb U878 ( .A(AD22I), .Y(n3437) );
    zor2b U879 ( .A(n3099), .B(n3323), .Y(n3091) );
    zivb U880 ( .A(n3091), .Y(n3100) );
    zmux21lb U881 ( .A(n3416), .B(n3432), .S(n2978), .Y(INTTHRESHOLD1414_1) );
    zivb U882 ( .A(AD17I), .Y(n3432) );
    zor2b U883 ( .A(n2982), .B(n3086), .Y(n_1613) );
    zivb U884 ( .A(n3077), .Y(n3080) );
    zivb U885 ( .A(n3323), .Y(n3329) );
    zmux21lb U886 ( .A(n3328), .B(n3439), .S(n3080), .Y(n3086) );
    zivb U887 ( .A(AD9I), .Y(n3439) );
    zmux21lb U888 ( .A(n3278), .B(n3428), .S(n2984), .Y(n_842) );
    zivb U889 ( .A(AD26I), .Y(n3428) );
    zmux21lb U890 ( .A(n3293), .B(n3438), .S(n2985), .Y(n_557) );
    zivb U891 ( .A(AD23I), .Y(n3438) );
    zmux21lb U892 ( .A(n3277), .B(n3427), .S(n2984), .Y(n_844) );
    zivb U893 ( .A(AD25I), .Y(n3427) );
    zivb U894 ( .A(AD15I), .Y(n3076) );
    zivb U895 ( .A(n3078), .Y(n3081) );
    zmux21lb U896 ( .A(n3313), .B(n3106), .S(n2987), .Y(n_1886) );
    zivb U897 ( .A(SUBIDWE), .Y(n3275) );
    zor2b U898 ( .A(n3040), .B(PORTCHG_S), .Y(USBSTS2) );
    zivb U899 ( .A(AD2I), .Y(n3106) );
    zor2b U900 ( .A(n3039), .B(ROLLOVER_S), .Y(USBSTS3) );
    zivb U901 ( .A(AD3I), .Y(n3109) );
    zor2b U902 ( .A(n3041), .B(HSERR_S), .Y(USBSTS4) );
    zivb U903 ( .A(AD4I), .Y(n3097) );
    zan2b U904 ( .A(n3074), .B(n3047), .Y(DBGPORT_R10G) );
    zivb U905 ( .A(n3374), .Y(n3074) );
    zivb U906 ( .A(PA4I), .Y(n3335) );
    zan2b U907 ( .A(n2989), .B(n3049), .Y(DBGPORT_R05G) );
    zan2b U908 ( .A(n3044), .B(n3045), .Y(DBGPORT_R04G) );
    zan2b U909 ( .A(n2995), .B(n3060), .Y(DBGPORT_R03G) );
    zivb U910 ( .A(n3273), .Y(n3060) );
    zor2b U911 ( .A(CBE3I_), .B(n3272), .Y(n3273) );
    zan2b U912 ( .A(n3044), .B(n3057), .Y(DBGPORT_R02G) );
    zan2b U913 ( .A(n3505), .B(n3049), .Y(DBGPORT_R01G) );
    zan2b U914 ( .A(n3044), .B(n3047), .Y(DBGPORT_R00G) );
    zivb U915 ( .A(n3368), .Y(n3044) );
    zivb U916 ( .A(PA7I), .Y(n3367) );
    zan2b U917 ( .A(UTM_RUN_T), .B(n3425), .Y(n3068) );
    zan2b U918 ( .A(n3046), .B(n3047), .Y(PSC_CBE0_H) );
    zan2b U919 ( .A(n2992), .B(n3049), .Y(PSC_CBE1_H) );
    zan2b U920 ( .A(n3046), .B(n3057), .Y(PSC_CBE2_H) );
    zivb U921 ( .A(n3379), .Y(n3046) );
    zan2b U922 ( .A(n3050), .B(n3055), .Y(PSC_CBE2_G) );
    zan2b U923 ( .A(n3058), .B(n3066), .Y(PSC_CBE0_F) );
    zan2b U924 ( .A(n3059), .B(n3049), .Y(PSC_CBE1_F) );
    zan2b U925 ( .A(n3058), .B(n3045), .Y(PSC_CBE0_E) );
    zan2b U926 ( .A(n3511), .B(n3049), .Y(PSC_CBE1_E) );
    zan2b U927 ( .A(n3005), .B(n3055), .Y(PSC_CBE2_E) );
    zor2b U928 ( .A(n3320), .B(n3381), .Y(n3384) );
    zan2b U929 ( .A(n3058), .B(n3047), .Y(PSC_CBE0_D) );
    zan2b U930 ( .A(n3063), .B(n3049), .Y(PSC_CBE1_D) );
    zor2b U931 ( .A(n3271), .B(n3381), .Y(n3385) );
    zan2b U932 ( .A(n3058), .B(n3057), .Y(PSC_CBE2_D) );
    zivb U933 ( .A(n3381), .Y(n3058) );
    zivb U934 ( .A(n3285), .Y(n3057) );
    zor2b U935 ( .A(n3271), .B(n3284), .Y(n3285) );
    zan2b U936 ( .A(n3507), .B(n3051), .Y(PSC_CBE0_C) );
    zivb U937 ( .A(n3309), .Y(n3051) );
    zor2b U938 ( .A(CBE0I_), .B(n3272), .Y(n3309) );
    zan2b U939 ( .A(n3053), .B(n3066), .Y(PSC_CBE0_B) );
    zivb U940 ( .A(n3310), .Y(n3066) );
    zor2b U941 ( .A(n3295), .B(n3309), .Y(n3310) );
    zan2b U942 ( .A(n3510), .B(n3049), .Y(PSC_CBE1_B) );
    zan2b U943 ( .A(n3053), .B(n3045), .Y(PSC_CBE0_A) );
    zivb U944 ( .A(n3332), .Y(n3045) );
    zor2b U945 ( .A(n3309), .B(n3320), .Y(n3332) );
    zan2b U946 ( .A(n3001), .B(n3049), .Y(PSC_CBE1_A) );
    zivb U947 ( .A(n3296), .Y(n3049) );
    zor2b U948 ( .A(CBE1I_), .B(n3272), .Y(n3296) );
    zan2b U949 ( .A(n3509), .B(n3055), .Y(PSC_CBE2_A) );
    zor2b U950 ( .A(n3320), .B(n3386), .Y(n3389) );
    zivb U951 ( .A(n3284), .Y(n3055) );
    zor2b U952 ( .A(CBE2I_), .B(n3272), .Y(n3284) );
    zivb U953 ( .A(REGW), .Y(n3272) );
    zan2b U954 ( .A(n3053), .B(n3047), .Y(CFG_CS) );
    zivb U955 ( .A(n3386), .Y(n3053) );
    zivb U956 ( .A(PA6I), .Y(n3378) );
    zivb U957 ( .A(n3366), .Y(n3047) );
    zor2b U958 ( .A(n3271), .B(n3309), .Y(n3366) );
    zivb U959 ( .A(n3424), .Y(HCHALT) );
    znd3b U960 ( .A(EHCI_IDLE), .B(n3425), .C(MAC_EOT), .Y(n3424) );
    zor2b U961 ( .A(n3070), .B(n3071), .Y(UINTOE_) );
    zivb U962 ( .A(UIRQACT), .Y(n3070) );
    zan2b U963 ( .A(n3072), .B(n3073), .Y(WR_ASYNCADDR) );
    zivb U964 ( .A(n3341), .Y(n3072) );
    zivb U965 ( .A(PA5I), .Y(n3340) );
    zivb U966 ( .A(n3295), .Y(n3073) );
    zor2b U967 ( .A(PA2I), .B(n3294), .Y(n3295) );
    zivb U968 ( .A(PA3I), .Y(n3294) );
    zan2b U969 ( .A(n2979), .B(n3061), .Y(WR_FRNUM) );
    zivb U970 ( .A(n3339), .Y(n3061) );
    zao22b U971 ( .A(HCCPARAMS_0), .B(n3450), .C(n3458), .D(USBINT_EN), .Y(
        n3111) );
    zao22b U972 ( .A(FRNUM_SYNC_0), .B(n2979), .C(PORTSC1[0]), .D(n3002), .Y(
        n3113) );
    zao22b U973 ( .A(DBGPORT_BUF1[2]), .B(n3447), .C(DBGPORT_ADDR[2]), .D(
        n3506), .Y(n3121) );
    zao22b U974 ( .A(PORTSC4[3]), .B(n2998), .C(PORTSC5[3]), .D(n3005), .Y(
        n3124) );
    zao22b U975 ( .A(DBGPORT_BUF1[3]), .B(n3447), .C(DBGPORT_ADDR[3]), .D(
        n3506), .Y(n3125) );
    zivb U976 ( .A(n3394), .Y(n3459) );
    zao22b U977 ( .A(HCCPARAMS_4), .B(n3450), .C(n3458), .D(HSERR_EN), .Y(
        n3128) );
    zivb U978 ( .A(n3393), .Y(n3458) );
    zao22b U979 ( .A(FRNUM_SYNC_4), .B(n2979), .C(PORTSC1[4]), .D(n3002), .Y(
        n3130) );
    zao2x4b U980 ( .A(INTDOORBELL), .B(n3452), .C(HCCPARAMS_6), .D(n3450), .E(
        HCSPARAMS_6), .F(n3451), .G(FRNUM_SYNC_6), .H(n2979), .Y(n3137) );
    zao22b U981 ( .A(DBGPORT_BUF1[6]), .B(n3447), .C(DBGPORT_ADDR[6]), .D(
        n3506), .Y(n3141) );
    zao2x4b U982 ( .A(n3452), .B(LIGHTRST), .C(HCCPARAMS_7), .D(n3450), .E(
        HCSPARAMS_7), .F(n3451), .G(FRNUM_SYNC_7), .H(n2979), .Y(n3143) );
    znd5b U983 ( .A(n3149), .B(n3150), .C(n3151), .D(n3152), .E(n3153), .Y(
        REGDOUT2[8]) );
    zaoi222b U984 ( .A(DBGPORT_BUF2[8]), .B(n3448), .C(DBGPORT_PID[8]), .D(
        n2989), .E(DBGPORT_SC[8]), .F(n3505), .Y(n3151) );
    zaoi22b U985 ( .A(DBGPORT_ADDR[8]), .B(n3506), .C(DBGPORT_BUF1[8]), .D(
        n3513), .Y(n3152) );
    znd5b U986 ( .A(n3154), .B(n3155), .C(n3156), .D(n3157), .E(n3158), .Y(
        REGDOUT2[9]) );
    zaoi222b U987 ( .A(DBGPORT_BUF2[9]), .B(n3514), .C(n3069), .D(DBGPORT_PID
        [9]), .E(n2996), .F(DBGPORT_SC[9]), .Y(n3156) );
    zaoi22b U988 ( .A(n3506), .B(DBGPORT_ADDR[9]), .C(DBGPORT_BUF1[9]), .D(
        n3447), .Y(n3157) );
    zaoi2x4b U989 ( .A(n2993), .B(PORTSC8[9]), .C(n3010), .D(PORTSC7[9]), .E(
        n3008), .F(PORTSC6[9]), .G(n3006), .H(PORTSC5[9]), .Y(n3158) );
    znd5b U990 ( .A(n3159), .B(n3160), .C(n3161), .D(n3162), .E(n3163), .Y(
        REGDOUT2[10]) );
    zaoi222b U991 ( .A(DBGPORT_BUF2[10]), .B(n3514), .C(DBGPORT_PID[10]), .D(
        n3069), .E(DBGPORT_SC[10]), .F(n2996), .Y(n3161) );
    znd5b U992 ( .A(n3164), .B(n3165), .C(n3166), .D(n3167), .E(n3168), .Y(
        REGDOUT2[11]) );
    zivb U993 ( .A(n3297), .Y(n3450) );
    zivb U994 ( .A(n3321), .Y(n3451) );
    zaoi222b U995 ( .A(DBGPORT_BUF2[11]), .B(n3448), .C(DBGPORT_PID[11]), .D(
        n2989), .E(DBGPORT_SC[11]), .F(n2996), .Y(n3166) );
    zaoi22b U996 ( .A(DBGPORT_ADDR[11]), .B(n3506), .C(DBGPORT_BUF1[11]), .D(
        n3513), .Y(n3167) );
    zao22b U997 ( .A(DBGPORT_BUF1[12]), .B(n3447), .C(DBGPORT_ADDR[12]), .D(
        n3506), .Y(n3171) );
    zoai2x4b U998 ( .A(n3266), .B(n3394), .C(n3321), .D(n3331), .E(n3396), .F(
        n3421), .G(n3297), .H(n3307), .Y(n3177) );
    zao22b U999 ( .A(DBGPORT_BUF1[14]), .B(n3447), .C(DBGPORT_ADDR[14]), .D(
        n3506), .Y(n3181) );
    zoai2x4b U1000 ( .A(n3268), .B(n3394), .C(n3321), .D(n3079), .E(n3396), 
        .F(n3420), .G(n3297), .H(n3308), .Y(n3183) );
    znd5b U1001 ( .A(n3189), .B(n3190), .C(n3191), .D(n3192), .E(n3193), .Y(
        REGDOUT2[16]) );
    zaoi222b U1002 ( .A(DBGPORT_BUF2[16]), .B(n3514), .C(DBGPORT_PID[16]), .D(
        n2990), .E(DBGPORT_SC[16]), .F(n3505), .Y(n3191) );
    znd5b U1003 ( .A(n3194), .B(n3195), .C(n3196), .D(n3197), .E(n3198), .Y(
        REGDOUT2[17]) );
    zaoi222b U1004 ( .A(DBGPORT_BUF2[17]), .B(n3448), .C(DBGPORT_PID[17]), .D(
        n2990), .E(DBGPORT_SC[17]), .F(n2996), .Y(n3196) );
    zaoi22b U1005 ( .A(DBGPORT_ADDR[17]), .B(n3506), .C(DBGPORT_BUF1[17]), .D(
        n3513), .Y(n3197) );
    znd5b U1006 ( .A(n3199), .B(n3200), .C(n3201), .D(n3202), .E(n3203), .Y(
        REGDOUT2[18]) );
    zaoi222b U1007 ( .A(DBGPORT_BUF2[18]), .B(n3514), .C(DBGPORT_PID[18]), .D(
        n2989), .E(DBGPORT_SC[18]), .F(n2996), .Y(n3201) );
    znd5b U1008 ( .A(n3204), .B(n3205), .C(n3206), .D(n3207), .E(n3208), .Y(
        REGDOUT2[19]) );
    zaoi222b U1009 ( .A(DBGPORT_BUF2[19]), .B(n3448), .C(DBGPORT_PID[19]), .D(
        n3069), .E(DBGPORT_SC[19]), .F(n2995), .Y(n3206) );
    zaoi22b U1010 ( .A(DBGPORT_ADDR[19]), .B(n3506), .C(DBGPORT_BUF1[19]), .D(
        n3513), .Y(n3207) );
    zoai2x4b U1011 ( .A(n3321), .B(n3370), .C(n3396), .D(n3411), .E(n3274), 
        .F(n3290), .G(n3391), .H(n3410), .Y(n3211) );
    zivb U1012 ( .A(EN_DBG_PORT), .Y(n3370) );
    znd5b U1013 ( .A(n3215), .B(n3216), .C(n3217), .D(n3218), .E(n3219), .Y(
        REGDOUT2[21]) );
    zaoi222b U1014 ( .A(DBGPORT_BUF2[21]), .B(n3514), .C(DBGPORT_PID[21]), .D(
        n2989), .E(DBGPORT_SC[21]), .F(n2995), .Y(n3217) );
    znd5b U1015 ( .A(n3220), .B(n3221), .C(n3222), .D(n3223), .E(n3224), .Y(
        REGDOUT2[22]) );
    zaoi222b U1016 ( .A(DBGPORT_BUF2[22]), .B(n3448), .C(DBGPORT_PID[22]), .D(
        n3069), .E(DBGPORT_SC[22]), .F(n3505), .Y(n3222) );
    zaoi22b U1017 ( .A(DBGPORT_ADDR[22]), .B(n3506), .C(DBGPORT_BUF1[22]), .D(
        n3513), .Y(n3223) );
    zivb U1018 ( .A(n3375), .Y(n3506) );
    zivb U1019 ( .A(n3373), .Y(n3513) );
    zivb U1020 ( .A(n3383), .Y(n3059) );
    znd5b U1021 ( .A(n3225), .B(n3226), .C(n3227), .D(n3228), .E(n3229), .Y(
        REGDOUT2[23]) );
    zivb U1022 ( .A(n3391), .Y(n3452) );
    zaoi222b U1023 ( .A(DBGPORT_BUF2[23]), .B(n3514), .C(DBGPORT_PID[23]), .D(
        n2990), .E(DBGPORT_SC[23]), .F(n2995), .Y(n3227) );
    zivb U1024 ( .A(n3373), .Y(n3447) );
    zivb U1025 ( .A(n3382), .Y(n3050) );
    zivb U1026 ( .A(n3387), .Y(n3507) );
    zivb U1027 ( .A(n3371), .Y(n3514) );
    zivb U1028 ( .A(n3388), .Y(n3510) );
    zivb U1029 ( .A(n3396), .Y(n3465) );
    zivb U1030 ( .A(n3274), .Y(n3460) );
    zivb U1031 ( .A(n3371), .Y(n3448) );
    zivb U1032 ( .A(INTASYNC), .Y(n3357) );
    zivb U1033 ( .A(ERRINT), .Y(n3355) );
    zivb U1034 ( .A(USBINT), .Y(n3358) );
    zdffqrb DBG_BUF_RG_reg_7 ( .CK(PCICLK), .D(RAFG), .R(HRST_), .Q(
        DBGPORT_R0FG) );
    zdffqrb DBG_BUF_RG_reg_6 ( .CK(PCICLK), .D(RAEG), .R(HRST_), .Q(
        DBGPORT_R0EG) );
    zdffqrb DBG_BUF_RG_reg_5 ( .CK(PCICLK), .D(RADG), .R(HRST_), .Q(
        DBGPORT_R0DG) );
    zdffqrb DBG_BUF_RG_reg_4 ( .CK(PCICLK), .D(RACG), .R(HRST_), .Q(
        DBGPORT_R0CG) );
    zdffqrb DBG_BUF_RG_reg_3 ( .CK(PCICLK), .D(RABG), .R(HRST_), .Q(
        DBGPORT_R0BG) );
    zdffqrb DBG_BUF_RG_reg_2 ( .CK(PCICLK), .D(RAAG), .R(HRST_), .Q(
        DBGPORT_R0AG) );
    zdffqrb DBG_BUF_RG_reg_1 ( .CK(PCICLK), .D(RA9G), .R(HRST_), .Q(
        DBGPORT_R09G) );
    zdffqrb DBG_BUF_RG_reg_0 ( .CK(PCICLK), .D(RA8G), .R(HRST_), .Q(
        DBGPORT_R08G) );
    zdffqsb ENUSB_reg_3 ( .CK(PCICLK), .D(ENUSB4), .S(HRST_), .Q(ENUSB_3) );
    zdffqsb ENUSB_reg_2 ( .CK(PCICLK), .D(ENUSB3), .S(HRST_), .Q(ENUSB_2) );
    zdffqsb ENUSB_reg_1 ( .CK(PCICLK), .D(ENUSB2), .S(HRST_), .Q(ENUSB_1) );
    zdffqsb ENUSB_reg_0 ( .CK(PCICLK), .D(ENUSB1), .S(HRST_), .Q(ENUSB_0) );
    zdffrb FRLSTSIZE_reg_1 ( .CK(PCICLK), .D(FRLSTSIZE1579_1), .R(n3525), .Q(
        FRLSTSIZE[1]), .QN(n3107) );
    zdffrb FRLSTSIZE_reg_0 ( .CK(PCICLK), .D(FRLSTSIZE1579_0), .R(CMDRST_), 
        .Q(FRLSTSIZE[0]), .QN(n3104) );
    zdffrb FLBASE_reg_31 ( .CK(PCICLK), .D(FLBASE2087_31), .R(n3525), .Q(
        FLBASE[31]), .QN(n3395) );
    zdffrb FLBASE_reg_30 ( .CK(PCICLK), .D(FLBASE2087_30), .R(n3524), .Q(
        FLBASE[30]), .QN(n3397) );
    zdffrb FLBASE_reg_29 ( .CK(PCICLK), .D(FLBASE2087_29), .R(CMDRST_), .Q(
        FLBASE[29]), .QN(n3398) );
    zdffrb FLBASE_reg_28 ( .CK(PCICLK), .D(FLBASE2087_28), .R(n3525), .Q(
        FLBASE[28]), .QN(n3399) );
    zdffrb FLBASE_reg_27 ( .CK(PCICLK), .D(FLBASE2087_27), .R(n3524), .Q(
        FLBASE[27]), .QN(n3400) );
    zdffrb FLBASE_reg_26 ( .CK(PCICLK), .D(FLBASE2087_26), .R(CMDRST_), .Q(
        FLBASE[26]), .QN(n3401) );
    zdffrb FLBASE_reg_25 ( .CK(PCICLK), .D(FLBASE2087_25), .R(n3525), .Q(
        FLBASE[25]), .QN(n3402) );
    zdffrb FLBASE_reg_24 ( .CK(PCICLK), .D(FLBASE2087_24), .R(n3524), .Q(
        FLBASE[24]), .QN(n3403) );
    zdffrb FLBASE_reg_23 ( .CK(PCICLK), .D(FLBASE2087_23), .R(CMDRST_), .Q(
        FLBASE[23]), .QN(n3405) );
    zdffrb FLBASE_reg_22 ( .CK(PCICLK), .D(FLBASE2087_22), .R(n3525), .Q(
        FLBASE[22]), .QN(n3407) );
    zdffrb FLBASE_reg_21 ( .CK(PCICLK), .D(FLBASE2087_21), .R(n3524), .Q(
        FLBASE[21]), .QN(n3409) );
    zdffrb FLBASE_reg_20 ( .CK(PCICLK), .D(FLBASE2087_20), .R(CMDRST_), .Q(
        FLBASE[20]), .QN(n3411) );
    zdffrb FLBASE_reg_19 ( .CK(PCICLK), .D(FLBASE2087_19), .R(n3525), .Q(
        FLBASE[19]), .QN(n3413) );
    zdffrb FLBASE_reg_18 ( .CK(PCICLK), .D(FLBASE2087_18), .R(n3524), .Q(
        FLBASE[18]), .QN(n3415) );
    zdffrb FLBASE_reg_17 ( .CK(PCICLK), .D(FLBASE2087_17), .R(CMDRST_), .Q(
        FLBASE[17]), .QN(n3417) );
    zdffrb FLBASE_reg_16 ( .CK(PCICLK), .D(FLBASE2087_16), .R(n3525), .Q(
        FLBASE[16]), .QN(n3419) );
    zdffrb FLBASE_reg_15 ( .CK(PCICLK), .D(FLBASE2087_15), .R(n3524), .Q(
        FLBASE[15]), .QN(n3420) );
    zdffrb FLBASE_reg_14 ( .CK(PCICLK), .D(FLBASE2087_14), .R(CMDRST_), .Q(
        FLBASE[14]), .QN(n3421) );
    zdffrb FLBASE_reg_13 ( .CK(PCICLK), .D(FLBASE2087_13), .R(n3525), .Q(
        FLBASE[13]), .QN(n3422) );
    zdffrb FLBASE_reg_12 ( .CK(PCICLK), .D(FLBASE2087_12), .R(n3524), .Q(
        FLBASE[12]), .QN(n3423) );
    zdffqb REGDOUT_reg_31 ( .CK(PCICLK), .D(REGDOUT2[31]), .Q(REGD31) );
    zdffqb REGDOUT_reg_30 ( .CK(PCICLK), .D(REGDOUT2[30]), .Q(REGD30) );
    zdffqb REGDOUT_reg_29 ( .CK(PCICLK), .D(REGDOUT2[29]), .Q(REGD29) );
    zdffqb REGDOUT_reg_28 ( .CK(PCICLK), .D(REGDOUT2[28]), .Q(REGD28) );
    zdffqb REGDOUT_reg_27 ( .CK(PCICLK), .D(REGDOUT2[27]), .Q(REGD27) );
    zdffqb REGDOUT_reg_26 ( .CK(PCICLK), .D(REGDOUT2[26]), .Q(REGD26) );
    zdffqb REGDOUT_reg_25 ( .CK(PCICLK), .D(REGDOUT2[25]), .Q(REGD25) );
    zdffqb REGDOUT_reg_24 ( .CK(PCICLK), .D(REGDOUT2[24]), .Q(REGD24) );
    zdffqb REGDOUT_reg_23 ( .CK(PCICLK), .D(REGDOUT2[23]), .Q(REGD23) );
    zdffqb REGDOUT_reg_22 ( .CK(PCICLK), .D(REGDOUT2[22]), .Q(REGD22) );
    zdffqb REGDOUT_reg_21 ( .CK(PCICLK), .D(REGDOUT2[21]), .Q(REGD21) );
    zdffqb REGDOUT_reg_20 ( .CK(PCICLK), .D(REGDOUT2[20]), .Q(REGD20) );
    zdffqb REGDOUT_reg_19 ( .CK(PCICLK), .D(REGDOUT2[19]), .Q(REGD19) );
    zdffqb REGDOUT_reg_18 ( .CK(PCICLK), .D(REGDOUT2[18]), .Q(REGD18) );
    zdffqb REGDOUT_reg_17 ( .CK(PCICLK), .D(REGDOUT2[17]), .Q(REGD17) );
    zdffqb REGDOUT_reg_16 ( .CK(PCICLK), .D(REGDOUT2[16]), .Q(REGD16) );
    zdffqb REGDOUT_reg_15 ( .CK(PCICLK), .D(REGDOUT2[15]), .Q(REGD15) );
    zdffqb REGDOUT_reg_14 ( .CK(PCICLK), .D(REGDOUT2[14]), .Q(REGD14) );
    zdffqb REGDOUT_reg_13 ( .CK(PCICLK), .D(REGDOUT2[13]), .Q(REGD13) );
    zdffqb REGDOUT_reg_12 ( .CK(PCICLK), .D(REGDOUT2[12]), .Q(REGD12) );
    zdffqb REGDOUT_reg_11 ( .CK(PCICLK), .D(REGDOUT2[11]), .Q(REGD11) );
    zdffqb REGDOUT_reg_10 ( .CK(PCICLK), .D(REGDOUT2[10]), .Q(REGD10) );
    zdffqb REGDOUT_reg_9 ( .CK(PCICLK), .D(REGDOUT2[9]), .Q(REGD9) );
    zdffqb REGDOUT_reg_8 ( .CK(PCICLK), .D(REGDOUT2[8]), .Q(REGD8) );
    zdffqb REGDOUT_reg_7 ( .CK(PCICLK), .D(REGDOUT2[7]), .Q(REGD7) );
    zdffqb REGDOUT_reg_6 ( .CK(PCICLK), .D(REGDOUT2[6]), .Q(REGD6) );
    zdffqb REGDOUT_reg_5 ( .CK(PCICLK), .D(REGDOUT2[5]), .Q(REGD5) );
    zdffqb REGDOUT_reg_4 ( .CK(PCICLK), .D(REGDOUT2[4]), .Q(REGD4) );
    zdffqb REGDOUT_reg_3 ( .CK(PCICLK), .D(REGDOUT2[3]), .Q(REGD3) );
    zdffqb REGDOUT_reg_2 ( .CK(PCICLK), .D(REGDOUT2[2]), .Q(REGD2) );
    zdffqb REGDOUT_reg_1 ( .CK(PCICLK), .D(REGDOUT2[1]), .Q(REGD1) );
    zdffqb REGDOUT_reg_0 ( .CK(PCICLK), .D(REGDOUT2[0]), .Q(REGD0) );
    zdffqrb HCRESET_2T_reg ( .CK(PCICLK), .D(n3522), .R(HRST_), .Q(HCRESET_2T)
         );
    zdffrb HSERR_EN_reg ( .CK(PCICLK), .D(HSERR_EN2004), .R(CMDRST_), .Q(
        HSERR_EN), .QN(n3360) );
    zdffrb HCIVERSION_reg_5 ( .CK(PCICLK), .D(n_561), .R(HRST_), .Q(
        HCIVERSION_5), .QN(n3291) );
    zdffrb HCIVERSION_reg2_12 ( .CK(PCICLK), .D(n_838), .R(HRST_), .Q(
        HCIVERSION_12), .QN(n3280) );
    zdffrb HCSPARAMS_reg_6 ( .CK(PCICLK), .D(n_1238), .R(HRST_), .Q(
        HCSPARAMS_6), .QN(n3094) );
    zdffsb INTTHRESHOLD_reg_3 ( .CK(PCICLK), .D(INTTHRESHOLD1414_3), .S(n3525), 
        .Q(INTTHRESHOLD[3]), .QN(n3412) );
    zdffrb HCCPARAMS_reg2_15 ( .CK(PCICLK), .D(n_2151), .R(HRST_), .QN(n3308)
         );
    zdffqrb RUN_reg ( .CK(PCICLK_FREE), .D(RUN1760), .R(n3524), .Q(RUN) );
    zivb U1035 ( .A(RUN), .Y(n3425) );
    zdffqrb LIGHTRST_2T_reg ( .CK(PCICLK), .D(n3521), .R(HRST_), .Q(
        LIGHTRST_2T) );
    zdffrb SMIOWN_EN_reg ( .CK(PCICLK), .D(SMIOWN_EN2314), .R(HRST_), .Q(
        USBLEGCTLSTS[13]), .QN(n3343) );
    zdffrb HCCPARAMS_reg_0 ( .CK(PCICLK), .D(n_1890), .R(HRST_), .Q(
        HCCPARAMS_0), .QN(n3311) );
    zdffqrb USMIACT_T_reg ( .CK(PCICLK), .D(USMIACT), .R(HRST_), .Q(USMIACT_T)
         );
    zdffqrb SMIONBAR_reg ( .CK(PCICLK), .D(SMIONBAR_NXT), .R(HRST_), .Q(
        USBLEGCTLSTS[31]) );
    zivb U1036 ( .A(USBLEGCTLSTS[31]), .Y(n3347) );
    zdffrb HCSPARAMS_reg2_10 ( .CK(PCICLK), .D(n_1611), .R(HRST_), .Q(
        HCSPARAMS_10), .QN(n3085) );
    zdffqrb PERIOD_EN_reg ( .CK(PCICLK), .D(PERIOD_EN1619), .R(n3525), .Q(
        PERIOD_EN) );
    zivb U1037 ( .A(PERIOD_EN), .Y(n3265) );
    zdffrb HCCPARAMS_reg_7 ( .CK(PCICLK), .D(n_1876), .R(HRST_), .Q(
        HCCPARAMS_7), .QN(n3318) );
    zdffrb HCCPARAMS_reg2_12 ( .CK(PCICLK), .D(n_2157), .R(HRST_), .QN(n3303)
         );
    zdffrb INTDOORBELL_reg ( .CK(PCICLK_FREE), .D(INTDOORBELL1489), .R(n3525), 
        .Q(INTDOORBELL), .QN(n3392) );
    zdffrb SMIONPCMD_EN_reg ( .CK(PCICLK), .D(SMIONPCMD_EN2320), .R(HRST_), 
        .Q(USBLEGCTLSTS[14]), .QN(n3345) );
    zdffrb HCIVERSION_reg2_15 ( .CK(PCICLK), .D(n_832), .R(HRST_), .Q(
        HCIVERSION_15), .QN(n3283) );
    zdffrb INTTHRESHOLD_reg_4 ( .CK(PCICLK), .D(INTTHRESHOLD1414_4), .R(n3524), 
        .Q(INTTHRESHOLD[4]), .QN(n3410) );
    zdffqrb HCSPARAMS_reg_1 ( .CK(PCICLK), .D(n_1248), .R(HRST_), .Q(
        HCSPARAMS_1) );
    zdffrb USBINT_EN_reg ( .CK(PCICLK), .D(USBINT_EN1980), .R(CMDRST_), .Q(
        USBINT_EN), .QN(n3359) );
    zdffrb HCIVERSION_reg_2 ( .CK(PCICLK), .D(n_567), .R(HRST_), .Q(
        HCIVERSION_2), .QN(n3288) );
    zdffqrb OSOWNS_reg ( .CK(PCICLK), .D(OSOWNS2125), .R(HRST_), .Q(USBLEGSUP
        [24]) );
    zivb U1038 ( .A(USBLEGSUP[24]), .Y(n3441) );
    zdffqrb UTM_RUN_T_reg ( .CK(PCICLK), .D(RUN), .R(HRST_), .Q(UTM_RUN_T) );
    zdffsb HCCPARAMS_reg2_13 ( .CK(PCICLK), .D(n_2155), .S(HRST_), .Q(
        HCCPARAMS_13), .QN(n3305) );
    zdffrb ROLLOVER_EN_reg ( .CK(PCICLK), .D(ROLLOVER_EN1998), .R(n3525), .Q(
        ROLLOVER_EN), .QN(n3362) );
    zdffsb HCCPARAMS_reg_6 ( .CK(PCICLK), .D(n_1878), .S(HRST_), .Q(
        HCCPARAMS_6), .QN(n3317) );
    zdffqrb USMIO_2T_reg ( .CK(PCICLK), .D(n3520), .R(HRST_), .Q(USMIO_2T) );
    zdffrb HCSPARAMS_reg2_11 ( .CK(PCICLK), .D(n_1609), .R(HRST_), .Q(
        HCSPARAMS_11), .QN(n3083) );
    zdffqrb ASYNC_STS_reg ( .CK(PCICLK_FREE), .D(val1876_1), .R(n3524), .Q(
        ASYNC_STS) );
    zivb U1039 ( .A(ASYNC_STS), .Y(n3268) );
    zdffqrb FRNUM_PCLK_LATCH_33_reg ( .CK(PCICLK_FREE), .D(FRNUM_PCLK_LATCH_66
        ), .R(HRST_), .Q(n_3593) );
    zdffrb HCIVERSION_reg_3 ( .CK(PCICLK), .D(n_565), .R(HRST_), .Q(
        HCIVERSION_3), .QN(n3289) );
    zdffqrb SMIOSOWNCHG_reg ( .CK(PCICLK), .D(SMIOSOWNCHG_NXT), .R(HRST_), .Q(
        USBLEGCTLSTS[29]) );
    zivb U1040 ( .A(USBLEGCTLSTS[29]), .Y(n3342) );
    zdffrb SMIUSBERR_EN_reg ( .CK(PCICLK), .D(SMIUSBERR_EN2395), .R(HRST_), 
        .Q(USBLEGCTLSTS[1]), .QN(n3356) );
    zdffrb SMIFROVER_EN_reg ( .CK(PCICLK), .D(SMIFROVER_EN2407), .R(HRST_), 
        .Q(USBLEGCTLSTS[3]), .QN(n3354) );
    zdffrb HCIVERSION_reg2_14 ( .CK(PCICLK), .D(n_834), .R(HRST_), .Q(
        HCIVERSION_14), .QN(n3282) );
    zdffrb INTTHRESHOLD_reg_5 ( .CK(PCICLK), .D(INTTHRESHOLD1414_5), .R(n3524), 
        .Q(INTTHRESHOLD[5]), .QN(n3408) );
    zdffrb HCSPARAMS_reg_0 ( .CK(PCICLK), .D(n_1250), .R(HRST_), .Q(
        HCSPARAMS_0), .QN(n3102) );
    zdffrb HCIVERSION_reg2_13 ( .CK(PCICLK), .D(n_836), .R(HRST_), .Q(
        HCIVERSION_13), .QN(n3281) );
    zdffqrb LIGHTRST_T_reg ( .CK(PCICLK), .D(n3519), .R(HRST_), .Q(LIGHTRST_T)
         );
    zdffrb HCSPARAMS_reg_7 ( .CK(PCICLK), .D(n_1236), .R(HRST_), .Q(
        HCSPARAMS_7), .QN(n3092) );
    zdffrb INTTHRESHOLD_reg_2 ( .CK(PCICLK), .D(INTTHRESHOLD1414_2), .R(
        CMDRST_), .Q(INTTHRESHOLD[2]), .QN(n3414) );
    zdffqrb SMIONPCMD_reg ( .CK(PCICLK), .D(SMIONPCMD_NXT), .R(HRST_), .Q(
        USBLEGCTLSTS[30]) );
    zivb U1041 ( .A(USBLEGCTLSTS[30]), .Y(n3365) );
    zdffqrb BIOSOWNS_reg ( .CK(PCICLK), .D(BIOSOWNS2162), .R(HRST_), .Q(
        USBLEGSUP[16]) );
    zdffrb HCIVERSION_reg_4 ( .CK(PCICLK), .D(n_563), .R(HRST_), .QN(n3290) );
    zdffqrb_ USMIO_3T_reg ( .CK(PCICLK), .D(USMIO_T), .R(HRST_), .Q(USMIO_3T)
         );
    zdffqrb INTASYNC_EN_reg ( .CK(PCICLK), .D(INTASYNC_EN2010), .R(n3525), .Q(
        INTASYNC_EN) );
    zivb U1042 ( .A(INTASYNC_EN), .Y(n3363) );
    zdffsb HCCPARAMS_reg_1 ( .CK(PCICLK), .D(n_1888), .S(HRST_), .QN(n3312) );
    zdffqrb USMIO_T_reg ( .CK(PCICLK), .D(USMIO_T2541), .R(HRST_), .Q(USMIO_T)
         );
    zdffsb HCCPARAMS_reg2_14 ( .CK(PCICLK), .D(n_2153), .S(HRST_), .QN(n3307)
         );
    zdffqrb HCRESET_reg ( .CK(PCICLK), .D(HCRESET1670), .R(HRST_), .Q(HCRESET)
         );
    zivb U1043 ( .A(HCRESET), .Y(n_12) );
    zdffsb HCIVERSION_reg2_8 ( .CK(PCICLK), .D(n_846), .S(HRST_), .Q(
        HCIVERSION_8), .QN(n3276) );
    zdffqrb ASYNC_EN_reg ( .CK(PCICLK), .D(ASYNC_EN1625), .R(CMDRST_), .Q(
        ASYNC_EN) );
    zivb U1044 ( .A(ASYNC_EN), .Y(n3267) );
    zdffrb USBSMI_EN_reg ( .CK(PCICLK), .D(USBSMI_EN2389), .R(HRST_), .Q(
        USBLEGCTLSTS[0]), .QN(n3344) );
    zdffrb HCIVERSION_reg_6 ( .CK(PCICLK), .D(n_559), .R(HRST_), .Q(
        HCIVERSION_6), .QN(n3292) );
    zdffrb HCSPARAMS_reg_5 ( .CK(PCICLK), .D(n_1240), .R(HRST_), .Q(
        HCSPARAMS_5), .QN(n3096) );
    zdffrb INTTHRESHOLD_reg_0 ( .CK(PCICLK), .D(INTTHRESHOLD1414_0), .R(n3525), 
        .Q(INTTHRESHOLD[0]), .QN(n3418) );
    zdffrb HCIVERSION_reg2_11 ( .CK(PCICLK), .D(n_840), .R(HRST_), .Q(
        HCIVERSION_11), .QN(n3279) );
    zdffrb HCSPARAMS_reg2_8 ( .CK(PCICLK), .D(n_1615), .R(HRST_), .Q(
        HCSPARAMS_8), .QN(n3088) );
    zdffrb HCCPARAMS_reg_3 ( .CK(PCICLK), .D(n_1884), .R(HRST_), .QN(n3314) );
    zdffqsb HCSPARAMS_reg2_14 ( .CK(PCICLK), .D(n_1603), .S(HRST_), .Q(
        HCSPARAMS_14) );
    zivb U1045 ( .A(HCSPARAMS_14), .Y(n3331) );
    zdffrb SMIPORTCHG_EN_reg ( .CK(PCICLK), .D(SMIPORTCHG_EN2401), .R(HRST_), 
        .Q(USBLEGCTLSTS[2]), .QN(n3350) );
    zdffrb PORTCHG_EN_reg ( .CK(PCICLK), .D(PORTCHG_EN1992), .R(n3524), .Q(
        PORTCHG_EN), .QN(n3361) );
    zdffqrb HCSPARAMS_reg2_13 ( .CK(PCICLK), .D(n_1605), .R(HRST_), .Q(
        HCSPARAMS_13) );
    zdffsb HCCPARAMS_reg_4 ( .CK(PCICLK), .D(n_1882), .S(HRST_), .Q(
        HCCPARAMS_4), .QN(n3315) );
    zdffrb HCCPARAMS_reg2_9 ( .CK(PCICLK), .D(n_2163), .R(HRST_), .Q(
        HCCPARAMS_9), .QN(n3299) );
    zdffsb HCCPARAMS_reg2_11 ( .CK(PCICLK), .D(n_2159), .S(HRST_), .Q(
        HCCPARAMS_11), .QN(n3301) );
    zdffqrb HCSPARAMS_reg_2 ( .CK(PCICLK), .D(n_1246), .R(HRST_), .Q(
        HCSPARAMS_2) );
    zivb U1046 ( .A(HCSPARAMS_2), .Y(n3333) );
    zdffrb INTTHRESHOLD_reg_7 ( .CK(PCICLK), .D(INTTHRESHOLD1414_7), .R(
        CMDRST_), .Q(INTTHRESHOLD[7]), .QN(n3404) );
    zdffqrb PERIOD_STS_reg ( .CK(PCICLK_FREE), .D(val1944_1), .R(n3524), .Q(
        PERIOD_STS) );
    zivb U1047 ( .A(PERIOD_STS), .Y(n3266) );
    zdffrb HCIVERSION_reg_1 ( .CK(PCICLK), .D(n_569), .R(HRST_), .Q(
        HCIVERSION_1), .QN(n3287) );
    zdffrb SMIONBAR_EN_reg ( .CK(PCICLK), .D(SMIONBAR_EN2326), .R(HRST_), .Q(
        USBLEGCTLSTS[15]), .QN(n3348) );
    zdffrb SMIASYNC_EN_reg ( .CK(PCICLK), .D(SMIASYNC_EN2419), .R(HRST_), .Q(
        USBLEGCTLSTS[5]), .QN(n3346) );
    zdffrb HCCPARAMS_reg2_8 ( .CK(PCICLK), .D(n_2165), .R(HRST_), .Q(
        HCCPARAMS_8), .QN(n3298) );
    zdffqrb LIGHTRST_reg ( .CK(PCICLK), .D(LIGHTRST1452), .R(HRST_), .Q(
        LIGHTRST) );
    zivb U1048 ( .A(LIGHTRST), .Y(n_14) );
    zdffrb HCCPARAMS_reg2_10 ( .CK(PCICLK), .D(n_2161), .R(HRST_), .Q(
        HCCPARAMS_10), .QN(n3300) );
    zdffsb HCCPARAMS_reg_5 ( .CK(PCICLK), .D(n_1880), .S(HRST_), .Q(
        HCCPARAMS_5), .QN(n3316) );
    zdffqrb HCSPARAMS_reg2_12 ( .CK(PCICLK), .D(n_1607), .R(HRST_), .Q(
        HCSPARAMS_12) );
    zivb U1049 ( .A(HCSPARAMS_12), .Y(n3330) );
    zdffrb HCIVERSION_reg_0 ( .CK(PCICLK), .D(n_571), .R(HRST_), .Q(
        HCIVERSION_0), .QN(n3286) );
    zdffrb ERRINT_EN_reg ( .CK(PCICLK), .D(ERRINT_EN1986), .R(n3525), .Q(
        ERRINT_EN), .QN(n3364) );
    zdffrb SMIHERR_EN_reg ( .CK(PCICLK), .D(SMIHERR_EN2413), .R(HRST_), .Q(
        USBLEGCTLSTS[4]), .QN(n3352) );
    zdffqsb HCSPARAMS_reg_3 ( .CK(PCICLK), .D(n_1244), .S(HRST_), .Q(
        HCSPARAMS_3) );
    zivb U1050 ( .A(HCSPARAMS_3), .Y(n3334) );
    zdffrb INTTHRESHOLD_reg_6 ( .CK(PCICLK), .D(INTTHRESHOLD1414_6), .R(n3524), 
        .Q(INTTHRESHOLD[6]), .QN(n3406) );
    zdffrb HCSPARAMS_reg_4 ( .CK(PCICLK), .D(n_1242), .R(HRST_), .Q(
        HCSPARAMS_4), .QN(n3098) );
    zdffrb INTTHRESHOLD_reg_1 ( .CK(PCICLK), .D(INTTHRESHOLD1414_1), .R(
        CMDRST_), .Q(INTTHRESHOLD[1]), .QN(n3416) );
    zdffsb HCSPARAMS_reg2_9 ( .CK(PCICLK), .D(n_1613), .S(HRST_), .Q(
        HCSPARAMS_9), .QN(n3328) );
    zdffrb HCIVERSION_reg2_10 ( .CK(PCICLK), .D(n_842), .R(HRST_), .Q(
        HCIVERSION_10), .QN(n3278) );
    zdffrb HCIVERSION_reg_7 ( .CK(PCICLK), .D(n_557), .R(HRST_), .Q(
        HCIVERSION_7), .QN(n3293) );
    zdffrb HCIVERSION_reg2_9 ( .CK(PCICLK), .D(n_844), .R(HRST_), .Q(
        HCIVERSION_9), .QN(n3277) );
    zdffrb HCSPARAMS_reg2_15 ( .CK(PCICLK), .D(n_1601), .R(HRST_), .QN(n3079)
         );
    zdffrb HCCPARAMS_reg_2 ( .CK(PCICLK), .D(n_1886), .R(HRST_), .QN(n3313) );
    zdffqrb HCRESET_T_reg ( .CK(PCICLK), .D(n3517), .R(HRST_), .Q(HCRESET_T)
         );
    zdffqrb sts2 ( .CK(PCICLK_FREE), .D(USBSTS2), .R(n3525), .Q(USBLEGCTLSTS
        [18]) );
    zivb U1051 ( .A(USBLEGCTLSTS[18]), .Y(n3349) );
    zdffqrb sts3 ( .CK(PCICLK_FREE), .D(USBSTS3), .R(CMDRST_), .Q(USBLEGCTLSTS
        [19]) );
    zivb U1052 ( .A(USBLEGCTLSTS[19]), .Y(n3353) );
    zdffqrb sts4 ( .CK(PCICLK_FREE), .D(USBSTS4), .R(n3524), .Q(USBLEGCTLSTS
        [20]) );
    zivb U1053 ( .A(USBLEGCTLSTS[20]), .Y(n3351) );
    znr2b U1054 ( .A(n3310), .B(n3338), .Y(n2977) );
    znr2b U1055 ( .A(n3285), .B(n3338), .Y(n2978) );
    znr2d U1056 ( .A(n3337), .B(n3338), .Y(n2979) );
    zoa21b U1057 ( .A(ENUSB2), .B(ENUSB3), .C(n3322), .Y(n2980) );
    znr2b U1058 ( .A(ENUSB4), .B(n3254), .Y(n2981) );
    znr2b U1059 ( .A(n3080), .B(n3329), .Y(n2982) );
    znr2b U1060 ( .A(n3329), .B(n3099), .Y(n2983) );
    znr3d U1061 ( .A(n3275), .B(n3274), .C(n3273), .Y(n2984) );
    znr3d U1062 ( .A(n3270), .B(n3275), .C(n3285), .Y(n2985) );
    znr3d U1063 ( .A(n3275), .B(n3297), .C(n3296), .Y(n2986) );
    znr3d U1064 ( .A(n3270), .B(n3275), .C(n3310), .Y(n2987) );
    ziv11b U1065 ( .A(n3376), .Y(n2989), .Z(n2988) );
    zivb U1066 ( .A(n2988), .Y(n2990) );
    zivb U1067 ( .A(n3376), .Y(n3069) );
    zor2b U1068 ( .A(n3320), .B(n3368), .Y(n3376) );
    ziv11b U1069 ( .A(n3380), .Y(n2992), .Z(n2991) );
    zivb U1070 ( .A(n2991), .Y(n2993) );
    zivb U1071 ( .A(n3380), .Y(n3067) );
    zor2b U1072 ( .A(n3271), .B(n3379), .Y(n3380) );
    ziv11b U1073 ( .A(n3377), .Y(n2995), .Z(n2994) );
    zivb U1074 ( .A(n2994), .Y(n2996) );
    zivb U1075 ( .A(n3377), .Y(n3505) );
    zor2b U1076 ( .A(n3271), .B(n3368), .Y(n3377) );
    ziv11b U1077 ( .A(n3385), .Y(n2998), .Z(n2997) );
    zivb U1078 ( .A(n2997), .Y(n2999) );
    zao22b U1079 ( .A(PORTSC4[13]), .B(n2998), .C(PORTSC5[13]), .D(n3006), .Y(
        n3174) );
    zao22b U1080 ( .A(PORTSC4[1]), .B(n3063), .C(PORTSC5[1]), .D(n3511), .Y(
        n3116) );
    zivb U1081 ( .A(n3385), .Y(n3063) );
    ziv11b U1082 ( .A(n3389), .Y(n3001), .Z(n3000) );
    zivb U1083 ( .A(n3000), .Y(n3002) );
    zao22b U1084 ( .A(PORTSC2[2]), .B(n3048), .C(PORTSC1[2]), .D(n3509), .Y(
        n3486) );
    zao22b U1085 ( .A(PORTSC2[12]), .B(n3048), .C(PORTSC1[12]), .D(n3509), .Y(
        n3494) );
    zao22b U1086 ( .A(PORTSC2[5]), .B(n3048), .C(PORTSC1[5]), .D(n3001), .Y(
        n3457) );
    zivb U1087 ( .A(n3389), .Y(n3509) );
    zivb U1088 ( .A(n3375), .Y(n3003) );
    zan2b U1089 ( .A(n3056), .B(n3049), .Y(DBGPORT_R11G) );
    zaoi22b U1090 ( .A(DBGPORT_ADDR[18]), .B(n3056), .C(DBGPORT_BUF1[18]), .D(
        n3447), .Y(n3202) );
    zaoi22b U1091 ( .A(DBGPORT_ADDR[16]), .B(n3056), .C(DBGPORT_BUF1[16]), .D(
        n3447), .Y(n3192) );
    zaoi22b U1092 ( .A(DBGPORT_ADDR[23]), .B(n3056), .C(DBGPORT_BUF1[23]), .D(
        n3447), .Y(n3228) );
    zaoi22b U1093 ( .A(DBGPORT_ADDR[10]), .B(n3056), .C(DBGPORT_BUF1[10]), .D(
        n3447), .Y(n3162) );
    zaoi22b U1094 ( .A(DBGPORT_ADDR[21]), .B(n3056), .C(DBGPORT_BUF1[21]), .D(
        n3447), .Y(n3218) );
    zao22b U1095 ( .A(DBGPORT_BUF1[7]), .B(n3513), .C(DBGPORT_ADDR[7]), .D(
        n3056), .Y(n3147) );
    zao22b U1096 ( .A(DBGPORT_BUF1[20]), .B(n3513), .C(DBGPORT_ADDR[20]), .D(
        n3056), .Y(n3213) );
    zao22b U1097 ( .A(DBGPORT_BUF1[15]), .B(n3513), .C(DBGPORT_ADDR[15]), .D(
        n3056), .Y(n3187) );
    zao22b U1098 ( .A(DBGPORT_BUF1[13]), .B(n3513), .C(DBGPORT_ADDR[13]), .D(
        n3056), .Y(n3175) );
    zao22b U1099 ( .A(DBGPORT_BUF1[1]), .B(n3513), .C(DBGPORT_ADDR[1]), .D(
        n3056), .Y(n3117) );
    zao22b U1100 ( .A(DBGPORT_BUF1[5]), .B(n3513), .C(DBGPORT_ADDR[5]), .D(
        n3056), .Y(n3135) );
    zor2b U1101 ( .A(n3271), .B(n3374), .Y(n3375) );
    zivb U1102 ( .A(n3375), .Y(n3056) );
    ziv11b U1103 ( .A(n3384), .Y(n3005), .Z(n3004) );
    zivb U1104 ( .A(n3004), .Y(n3006) );
    zao22b U1105 ( .A(PORTSC4[5]), .B(n2998), .C(PORTSC5[5]), .D(n3006), .Y(
        n3134) );
    zao22b U1106 ( .A(PORTSC4[12]), .B(n3063), .C(PORTSC5[12]), .D(n3006), .Y(
        n3170) );
    zao22b U1107 ( .A(PORTSC4[2]), .B(n2999), .C(PORTSC5[2]), .D(n3511), .Y(
        n3120) );
    zivb U1108 ( .A(n3384), .Y(n3511) );
    zivb U1109 ( .A(n3388), .Y(n3007) );
    zan2b U1110 ( .A(n3007), .B(n3055), .Y(PSC_CBE2_B) );
    zaoi2x4b U1111 ( .A(n2998), .B(PORTSC4[9]), .C(n3009), .D(PORTSC3[9]), .E(
        n3007), .F(PORTSC2[9]), .G(n3509), .H(PORTSC1[9]), .Y(n3155) );
    zaoi2x4b U1112 ( .A(PORTSC4[23]), .B(n2999), .C(PORTSC3[23]), .D(n3507), 
        .E(PORTSC2[23]), .F(n3510), .G(PORTSC1[23]), .H(n3001), .Y(n3226) );
    zaoi2x4b U1113 ( .A(PORTSC4[16]), .B(n3063), .C(PORTSC3[16]), .D(n3507), 
        .E(PORTSC2[16]), .F(n3510), .G(PORTSC1[16]), .H(n3509), .Y(n3190) );
    zaoi2x4b U1114 ( .A(PORTSC4[18]), .B(n2998), .C(PORTSC3[18]), .D(n3507), 
        .E(PORTSC2[18]), .F(n3007), .G(PORTSC1[18]), .H(n3001), .Y(n3200) );
    zaoi2x4b U1115 ( .A(PORTSC4[21]), .B(n2999), .C(PORTSC3[21]), .D(n3009), 
        .E(PORTSC2[21]), .F(n3007), .G(PORTSC1[21]), .H(n3002), .Y(n3216) );
    zaoi2x4b U1116 ( .A(PORTSC4[10]), .B(n3063), .C(PORTSC3[10]), .D(n3009), 
        .E(PORTSC2[10]), .F(n3510), .G(PORTSC1[10]), .H(n3509), .Y(n3160) );
    zao2x4b U1117 ( .A(PORTSC2[30]), .B(n3510), .C(PORTSC3[30]), .D(n3507), 
        .E(PORTSC4[30]), .F(n3063), .G(PORTSC5[30]), .H(n3005), .Y(n3248) );
    zao2x4b U1118 ( .A(PORTSC2[28]), .B(n3007), .C(PORTSC3[28]), .D(n3507), 
        .E(PORTSC4[28]), .F(n2998), .G(PORTSC5[28]), .H(n3511), .Y(n3242) );
    zao2x4b U1119 ( .A(PORTSC2[26]), .B(n3510), .C(PORTSC3[26]), .D(n3009), 
        .E(PORTSC4[26]), .F(n2999), .G(PORTSC5[26]), .H(n3006), .Y(n3236) );
    zao2x4b U1120 ( .A(PORTSC2[24]), .B(n3007), .C(PORTSC3[24]), .D(n3009), 
        .E(PORTSC4[24]), .F(n3063), .G(PORTSC5[24]), .H(n3005), .Y(n3230) );
    zao22b U1121 ( .A(PORTSC2[13]), .B(n3048), .C(PORTSC1[13]), .D(n3001), .Y(
        n3490) );
    zao22b U1122 ( .A(PORTSC2[3]), .B(n3048), .C(PORTSC1[3]), .D(n3001), .Y(
        n3470) );
    zao22b U1123 ( .A(PORTSC2[1]), .B(n3048), .C(PORTSC1[1]), .D(n3509), .Y(
        n3498) );
    zor2b U1124 ( .A(n3295), .B(n3386), .Y(n3388) );
    zivb U1125 ( .A(n3388), .Y(n3048) );
    zivb U1126 ( .A(n3383), .Y(n3008) );
    zan2b U1127 ( .A(n3008), .B(n3055), .Y(PSC_CBE2_F) );
    zaoi2x4b U1128 ( .A(PORTSC8[18]), .B(n2993), .C(PORTSC7[18]), .D(n3050), 
        .E(PORTSC6[18]), .F(n3059), .G(PORTSC5[18]), .H(n3511), .Y(n3203) );
    zaoi2x4b U1129 ( .A(PORTSC8[16]), .B(n2992), .C(PORTSC7[16]), .D(n3050), 
        .E(PORTSC6[16]), .F(n3059), .G(PORTSC5[16]), .H(n3511), .Y(n3193) );
    zaoi2x4b U1130 ( .A(PORTSC8[23]), .B(n2992), .C(PORTSC7[23]), .D(n3050), 
        .E(PORTSC6[23]), .F(n3008), .G(PORTSC5[23]), .H(n3006), .Y(n3229) );
    zaoi2x4b U1131 ( .A(PORTSC8[10]), .B(n2993), .C(PORTSC7[10]), .D(n3010), 
        .E(PORTSC6[10]), .F(n3008), .G(PORTSC5[10]), .H(n3511), .Y(n3163) );
    zaoi2x4b U1132 ( .A(PORTSC8[21]), .B(n3067), .C(PORTSC7[21]), .D(n3010), 
        .E(PORTSC6[21]), .F(n3059), .G(PORTSC5[21]), .H(n3006), .Y(n3219) );
    zao2x4b U1133 ( .A(PORTSC5[20]), .B(n3006), .C(PORTSC6[20]), .D(n3008), 
        .E(PORTSC7[20]), .F(n3050), .G(PORTSC8[20]), .H(n2992), .Y(n3212) );
    zao2x4b U1134 ( .A(PORTSC5[14]), .B(n3006), .C(PORTSC6[14]), .D(n3059), 
        .E(PORTSC7[14]), .F(n3050), .G(PORTSC8[14]), .H(n3067), .Y(n3180) );
    zao2x4b U1135 ( .A(PORTSC5[7]), .B(n3006), .C(PORTSC6[7]), .D(n3059), .E(
        PORTSC7[7]), .F(n3010), .G(PORTSC8[7]), .H(n2993), .Y(n3146) );
    zao2x4b U1136 ( .A(PORTSC6[29]), .B(n3008), .C(PORTSC7[29]), .D(n3050), 
        .E(PORTSC8[29]), .F(n3067), .G(DBGPORT_SC[29]), .H(n2996), .Y(n3473)
         );
    zao2x4b U1137 ( .A(PORTSC6[31]), .B(n3059), .C(PORTSC7[31]), .D(n3050), 
        .E(PORTSC8[31]), .F(n2992), .G(DBGPORT_SC[31]), .H(n3505), .Y(n3464)
         );
    zao2x4b U1138 ( .A(PORTSC6[27]), .B(n3008), .C(PORTSC7[27]), .D(n3010), 
        .E(PORTSC8[27]), .F(n2993), .G(DBGPORT_SC[27]), .H(n3505), .Y(n3477)
         );
    zao2x4b U1139 ( .A(PORTSC6[25]), .B(n3059), .C(PORTSC7[25]), .D(n3010), 
        .E(PORTSC8[25]), .F(n2993), .G(DBGPORT_SC[25]), .H(n2995), .Y(n3481)
         );
    zor2b U1140 ( .A(n3295), .B(n3381), .Y(n3383) );
    zivb U1141 ( .A(n3383), .Y(n3512) );
    zivb U1142 ( .A(n3387), .Y(n3009) );
    zan2b U1143 ( .A(n3009), .B(n3055), .Y(PSC_CBE2_C) );
    zan2b U1144 ( .A(n3009), .B(n3049), .Y(PSC_CBE1_C) );
    zaoi2x4b U1145 ( .A(PORTSC4[8]), .B(n3063), .C(PORTSC3[8]), .D(n3507), .E(
        PORTSC2[8]), .F(n3007), .G(PORTSC1[8]), .H(n3002), .Y(n3150) );
    zaoi2x4b U1146 ( .A(PORTSC4[17]), .B(n2998), .C(PORTSC3[17]), .D(n3009), 
        .E(PORTSC2[17]), .F(n3510), .G(PORTSC1[17]), .H(n3509), .Y(n3195) );
    zaoi2x4b U1147 ( .A(PORTSC4[22]), .B(n2999), .C(PORTSC3[22]), .D(n3009), 
        .E(PORTSC2[22]), .F(n3007), .G(PORTSC1[22]), .H(n3001), .Y(n3221) );
    zaoi2x4b U1148 ( .A(PORTSC4[19]), .B(n2998), .C(PORTSC3[19]), .D(n3507), 
        .E(PORTSC2[19]), .F(n3510), .G(PORTSC1[19]), .H(n3001), .Y(n3205) );
    zaoi2x4b U1149 ( .A(PORTSC4[11]), .B(n2999), .C(PORTSC3[11]), .D(n3507), 
        .E(PORTSC2[11]), .F(n3510), .G(PORTSC1[11]), .H(n3002), .Y(n3165) );
    zao2x4b U1150 ( .A(PORTSC2[31]), .B(n3510), .C(PORTSC3[31]), .D(n3009), 
        .E(PORTSC4[31]), .F(n3063), .G(PORTSC5[31]), .H(n3006), .Y(n3251) );
    zao2x4b U1151 ( .A(PORTSC2[25]), .B(n3007), .C(PORTSC3[25]), .D(n3507), 
        .E(PORTSC4[25]), .F(n2998), .G(PORTSC5[25]), .H(n3005), .Y(n3233) );
    zao2x4b U1152 ( .A(PORTSC2[29]), .B(n3007), .C(PORTSC3[29]), .D(n3507), 
        .E(PORTSC4[29]), .F(n2999), .G(PORTSC5[29]), .H(n3511), .Y(n3245) );
    zao2x4b U1153 ( .A(PORTSC2[27]), .B(n3007), .C(PORTSC3[27]), .D(n3009), 
        .E(PORTSC4[27]), .F(n2999), .G(PORTSC5[27]), .H(n3005), .Y(n3239) );
    zivb U1154 ( .A(n3387), .Y(n3062) );
    zor2b U1155 ( .A(n3337), .B(n3386), .Y(n3387) );
    zivb U1156 ( .A(n3382), .Y(n3010) );
    zan2b U1157 ( .A(n3010), .B(n3049), .Y(PSC_CBE1_G) );
    zan2b U1158 ( .A(n3010), .B(n3051), .Y(PSC_CBE0_G) );
    zaoi2x4b U1159 ( .A(PORTSC8[19]), .B(n2992), .C(PORTSC7[19]), .D(n3010), 
        .E(PORTSC6[19]), .F(n3059), .G(PORTSC5[19]), .H(n3005), .Y(n3208) );
    zaoi2x4b U1160 ( .A(PORTSC8[22]), .B(n3067), .C(PORTSC7[22]), .D(n3050), 
        .E(PORTSC6[22]), .F(n3059), .G(PORTSC5[22]), .H(n3511), .Y(n3224) );
    zaoi2x4b U1161 ( .A(PORTSC8[17]), .B(n2993), .C(PORTSC7[17]), .D(n3050), 
        .E(PORTSC6[17]), .F(n3008), .G(PORTSC5[17]), .H(n3511), .Y(n3198) );
    zaoi2x4b U1162 ( .A(PORTSC8[11]), .B(n2992), .C(PORTSC7[11]), .D(n3050), 
        .E(PORTSC6[11]), .F(n3008), .G(PORTSC5[11]), .H(n3005), .Y(n3168) );
    zaoi2x4b U1163 ( .A(PORTSC8[8]), .B(n3067), .C(PORTSC7[8]), .D(n3010), .E(
        PORTSC6[8]), .F(n3008), .G(PORTSC5[8]), .H(n3006), .Y(n3153) );
    zao2x4b U1164 ( .A(PORTSC5[6]), .B(n3006), .C(PORTSC6[6]), .D(n3008), .E(
        PORTSC7[6]), .F(n3050), .G(PORTSC8[6]), .H(n3067), .Y(n3140) );
    zao2x4b U1165 ( .A(PORTSC5[15]), .B(n3511), .C(PORTSC6[15]), .D(n3059), 
        .E(PORTSC7[15]), .F(n3010), .G(PORTSC8[15]), .H(n2993), .Y(n3186) );
    zao2x4b U1166 ( .A(PORTSC6[30]), .B(n3008), .C(PORTSC7[30]), .D(n3508), 
        .E(PORTSC8[30]), .F(n2992), .G(DBGPORT_SC[30]), .H(n2996), .Y(n3467)
         );
    zao2x4b U1167 ( .A(PORTSC6[28]), .B(n3008), .C(PORTSC7[28]), .D(n3050), 
        .E(PORTSC8[28]), .F(n2992), .G(DBGPORT_SC[28]), .H(n3505), .Y(n3475)
         );
    zao2x4b U1168 ( .A(PORTSC6[24]), .B(n3059), .C(PORTSC7[24]), .D(n3010), 
        .E(PORTSC8[24]), .F(n3067), .G(DBGPORT_SC[24]), .H(n2995), .Y(n3483)
         );
    zao2x4b U1169 ( .A(PORTSC6[26]), .B(n3059), .C(PORTSC7[26]), .D(n3050), 
        .E(PORTSC8[26]), .F(n3067), .G(DBGPORT_SC[26]), .H(n2995), .Y(n3479)
         );
    zao22b U1170 ( .A(PORTSC8[0]), .B(n3067), .C(PORTSC7[0]), .D(n3508), .Y(
        n3502) );
    zan2b U1171 ( .A(PORTSC7[4]), .B(n3508), .Y(n3263) );
    zor2b U1172 ( .A(n3337), .B(n3381), .Y(n3382) );
    zivb U1173 ( .A(n3382), .Y(n3508) );
    zivb U1174 ( .A(n3504), .Y(n3011) );
    zmux21lb U1175 ( .A(n3399), .B(n3430), .S(n3445), .Y(FLBASE2087_28) );
    zmux21lb U1176 ( .A(n3400), .B(n3429), .S(n3445), .Y(FLBASE2087_27) );
    zmux21lb U1177 ( .A(n3398), .B(n3257), .S(n3011), .Y(FLBASE2087_29) );
    zmux21lb U1178 ( .A(n3395), .B(n3260), .S(n3445), .Y(FLBASE2087_31) );
    zmux21lb U1179 ( .A(n3397), .B(n3262), .S(n3011), .Y(FLBASE2087_30) );
    zmux21lb U1180 ( .A(n3402), .B(n3427), .S(n3011), .Y(FLBASE2087_25) );
    zmux21lb U1181 ( .A(n3401), .B(n3428), .S(n3011), .Y(FLBASE2087_26) );
    zmux21lb U1182 ( .A(n3409), .B(n3436), .S(n3445), .Y(FLBASE2087_21) );
    zmux21lb U1183 ( .A(n3415), .B(n3433), .S(n3445), .Y(FLBASE2087_18) );
    zmux21lb U1184 ( .A(n3405), .B(n3438), .S(n3445), .Y(FLBASE2087_23) );
    zmux21lb U1185 ( .A(n3413), .B(n3434), .S(n3445), .Y(FLBASE2087_19) );
    zmux21lb U1186 ( .A(n3417), .B(n3432), .S(n3445), .Y(FLBASE2087_17) );
    zmux21lb U1187 ( .A(n3407), .B(n3437), .S(n3445), .Y(FLBASE2087_22) );
    zmux21lb U1188 ( .A(n3422), .B(n3304), .S(n3445), .Y(FLBASE2087_13) );
    zmux21lb U1189 ( .A(n3419), .B(n3431), .S(n3445), .Y(FLBASE2087_16) );
    zmux21lb U1190 ( .A(n3403), .B(n3426), .S(n3445), .Y(FLBASE2087_24) );
    zmux21lb U1191 ( .A(n3421), .B(n3306), .S(n3445), .Y(FLBASE2087_14) );
    zmux21lb U1192 ( .A(n3420), .B(n3076), .S(n3445), .Y(FLBASE2087_15) );
    zmux21lb U1193 ( .A(n3423), .B(n3302), .S(n3445), .Y(FLBASE2087_12) );
    zmux21lb U1194 ( .A(n3411), .B(n3435), .S(n3445), .Y(FLBASE2087_20) );
    zor2b U1195 ( .A(n3320), .B(n3341), .Y(n3504) );
    zivb U1196 ( .A(n3390), .Y(n3012) );
    zaoi2x4b U1197 ( .A(n3012), .B(ASYNCLISTADDR[9]), .C(FRNUM_SYNC_9), .D(
        n2979), .E(HCCPARAMS_9), .F(n3450), .G(HCSPARAMS_9), .H(n3451), .Y(
        n3154) );
    zaoi2x4b U1198 ( .A(ASYNCLISTADDR[21]), .B(n3012), .C(INTTHRESHOLD[5]), 
        .D(n3452), .E(HCIVERSION_5), .F(n3460), .G(FLBASE[21]), .H(n3465), .Y(
        n3215) );
    zaoi2x4b U1199 ( .A(ASYNCLISTADDR[16]), .B(n3012), .C(INTTHRESHOLD[0]), 
        .D(n3452), .E(HCIVERSION_0), .F(n3460), .G(FLBASE[16]), .H(n3465), .Y(
        n3189) );
    zaoi2x4b U1200 ( .A(ASYNCLISTADDR[22]), .B(n3012), .C(INTTHRESHOLD[6]), 
        .D(n3452), .E(HCIVERSION_6), .F(n3460), .G(FLBASE[22]), .H(n3465), .Y(
        n3220) );
    zaoi2x4b U1201 ( .A(ASYNCLISTADDR[19]), .B(n3012), .C(INTTHRESHOLD[3]), 
        .D(n3452), .E(HCIVERSION_3), .F(n3460), .G(FLBASE[19]), .H(n3465), .Y(
        n3204) );
    zaoi2x4b U1202 ( .A(ASYNCLISTADDR[18]), .B(n3012), .C(INTTHRESHOLD[2]), 
        .D(n3452), .E(HCIVERSION_2), .F(n3460), .G(FLBASE[18]), .H(n3465), .Y(
        n3199) );
    zaoi2x4b U1203 ( .A(ASYNCLISTADDR[8]), .B(n3012), .C(FRNUM_SYNC_8), .D(
        n2979), .E(HCCPARAMS_8), .F(n3450), .G(HCSPARAMS_8), .H(n3451), .Y(
        n3149) );
    zaoi2x4b U1204 ( .A(ASYNCLISTADDR[17]), .B(n3012), .C(INTTHRESHOLD[1]), 
        .D(n3452), .E(HCIVERSION_1), .F(n3460), .G(FLBASE[17]), .H(n3465), .Y(
        n3194) );
    zaoi2x4b U1205 ( .A(ASYNCLISTADDR[10]), .B(n3012), .C(FRNUM_SYNC_10), .D(
        n2979), .E(HCCPARAMS_10), .F(n3450), .G(HCSPARAMS_10), .H(n3451), .Y(
        n3159) );
    zaoi2x4b U1206 ( .A(ASYNCLISTADDR[11]), .B(n3012), .C(FRNUM_SYNC_11), .D(
        n2979), .E(HCCPARAMS_11), .F(n3450), .G(HCSPARAMS_11), .H(n3451), .Y(
        n3164) );
    zaoi2x4b U1207 ( .A(ASYNCLISTADDR[23]), .B(n3012), .C(INTTHRESHOLD[7]), 
        .D(n3452), .E(HCIVERSION_7), .F(n3460), .G(FLBASE[23]), .H(n3465), .Y(
        n3225) );
    zao2x4b U1208 ( .A(n3465), .B(FLBASE[31]), .C(HCIVERSION_15), .D(n3460), 
        .E(ASYNCLISTADDR[31]), .F(n3012), .G(PORTSC1[31]), .H(n3001), .Y(n3252
        ) );
    zao2x4b U1209 ( .A(FLBASE[24]), .B(n3465), .C(HCIVERSION_8), .D(n3460), 
        .E(ASYNCLISTADDR[24]), .F(n3449), .G(PORTSC1[24]), .H(n3509), .Y(n3231
        ) );
    zao2x4b U1210 ( .A(FLBASE[26]), .B(n3465), .C(HCIVERSION_10), .D(n3460), 
        .E(ASYNCLISTADDR[26]), .F(n3449), .G(PORTSC1[26]), .H(n3002), .Y(n3237
        ) );
    zao2x4b U1211 ( .A(FLBASE[30]), .B(n3465), .C(HCIVERSION_14), .D(n3460), 
        .E(ASYNCLISTADDR[30]), .F(n3449), .G(PORTSC1[30]), .H(n3002), .Y(n3249
        ) );
    zao2x4b U1212 ( .A(FLBASE[28]), .B(n3465), .C(HCIVERSION_12), .D(n3460), 
        .E(ASYNCLISTADDR[28]), .F(n3449), .G(PORTSC1[28]), .H(n3002), .Y(n3243
        ) );
    zao2x4b U1213 ( .A(FLBASE[25]), .B(n3465), .C(HCIVERSION_9), .D(n3460), 
        .E(ASYNCLISTADDR[25]), .F(n3449), .G(PORTSC1[25]), .H(n3509), .Y(n3234
        ) );
    zao2x4b U1214 ( .A(FLBASE[29]), .B(n3465), .C(HCIVERSION_13), .D(n3460), 
        .E(ASYNCLISTADDR[29]), .F(n3449), .G(PORTSC1[29]), .H(n3002), .Y(n3246
        ) );
    zao2x4b U1215 ( .A(FLBASE[27]), .B(n3465), .C(HCIVERSION_11), .D(n3460), 
        .E(ASYNCLISTADDR[27]), .F(n3449), .G(PORTSC1[27]), .H(n3001), .Y(n3240
        ) );
    zao22b U1216 ( .A(ASYNCLISTADDR[20]), .B(n3449), .C(PORTSC1[20]), .D(n3002
        ), .Y(n3210) );
    zao22b U1217 ( .A(ASYNCLISTADDR[6]), .B(n3449), .C(PORTSC1[6]), .D(n3509), 
        .Y(n3138) );
    zao22b U1218 ( .A(ASYNCLISTADDR[15]), .B(n3449), .C(PORTSC1[15]), .D(n3001
        ), .Y(n3184) );
    zao22b U1219 ( .A(ASYNCLISTADDR[14]), .B(n3449), .C(PORTSC1[14]), .D(n3002
        ), .Y(n3178) );
    zao22b U1220 ( .A(ASYNCLISTADDR[7]), .B(n3449), .C(PORTSC1[7]), .D(n3002), 
        .Y(n3144) );
    zivb U1221 ( .A(n3390), .Y(n3449) );
    zbfb U1222 ( .A(INTASYNC), .Y(USBLEGCTLSTS[21]) );
    zdffqrb sts5 ( .CK(PCICLK_FREE), .D(USBSTS5), .R(n3525), .Q(INTASYNC) );
    zbfb U1223 ( .A(ERRINT), .Y(USBLEGCTLSTS[17]) );
    zdffqrb sts1 ( .CK(PCICLK_FREE), .D(USBSTS1), .R(CMDRST_), .Q(ERRINT) );
    zbfb U1224 ( .A(USBINT), .Y(USBLEGCTLSTS[16]) );
    zdffqrb sts0 ( .CK(PCICLK_FREE), .D(USBSTS0), .R(n3524), .Q(USBINT) );
    zdffb FRNUM_SYNC_reg_13 ( .CK(PCICLK_FREE), .D(n3016), .Q(FRNUM_SYNC_13)
         );
    zdffb FRNUM_SYNC_reg_12 ( .CK(PCICLK_FREE), .D(n3017), .Q(FRNUM_SYNC_12)
         );
    zdffb FRNUM_SYNC_reg_11 ( .CK(PCICLK_FREE), .D(n3018), .Q(FRNUM_SYNC_11)
         );
    zdffb FRNUM_SYNC_reg_10 ( .CK(PCICLK_FREE), .D(n3019), .Q(FRNUM_SYNC_10)
         );
    zdffb FRNUM_SYNC_reg_9 ( .CK(PCICLK_FREE), .D(n3020), .Q(FRNUM_SYNC_9) );
    zdffb FRNUM_SYNC_reg_8 ( .CK(PCICLK_FREE), .D(n3021), .Q(FRNUM_SYNC_8) );
    zdffb FRNUM_SYNC_reg_7 ( .CK(PCICLK_FREE), .D(n3022), .Q(FRNUM_SYNC_7) );
    zdffb FRNUM_SYNC_reg_6 ( .CK(PCICLK_FREE), .D(n3023), .Q(FRNUM_SYNC_6) );
    zdffb FRNUM_SYNC_reg_5 ( .CK(PCICLK_FREE), .D(n3024), .Q(FRNUM_SYNC_5) );
    zdffb FRNUM_SYNC_reg_4 ( .CK(PCICLK_FREE), .D(n3025), .Q(FRNUM_SYNC_4) );
    zdffb FRNUM_SYNC_reg_3 ( .CK(PCICLK_FREE), .D(n3026), .Q(FRNUM_SYNC_3) );
    zdffb FRNUM_SYNC_reg_2 ( .CK(PCICLK_FREE), .D(n3027), .Q(FRNUM_SYNC_2) );
    zdffb FRNUM_SYNC_reg_1 ( .CK(PCICLK_FREE), .D(n3028), .Q(FRNUM_SYNC_1) );
    zdffb FRNUM_SYNC_reg_0 ( .CK(PCICLK_FREE), .D(n3029), .Q(FRNUM_SYNC_0) );
    zor4b U1225 ( .A(n3030), .B(n3031), .C(n3032), .D(n3033), .Y(USMIACT) );
    zor3b U1226 ( .A(USMIO_2T), .B(USMIO_3T), .C(USMIO_T), .Y(USMIO) );
    zao211b U1227 ( .A(INTASYNC_EN), .B(ASYNCINT), .C(n3064), .D(n3065), .Y(
        UIRQACT) );
    zinr2b U1228 ( .A(n3068), .B(DIS_SOF_RUN), .Y(UTM_RUN) );
    zoai22d U1229 ( .A(n3076), .B(n3077), .C(n3078), .D(n3079), .Y(n_1601) );
    zao222b U1230 ( .A(n3080), .B(AD14I), .C(n2982), .D(ENUSB4), .E(
        HCSPARAMS_14), .F(n3081), .Y(n_1603) );
    zao222b U1231 ( .A(n3080), .B(AD13I), .C(n2980), .D(n2982), .E(
        HCSPARAMS_13), .F(n3081), .Y(n_1605) );
    zao222b U1232 ( .A(n3080), .B(AD12I), .C(n2981), .D(n2982), .E(
        HCSPARAMS_12), .F(n3081), .Y(n_1607) );
    zoai22d U1233 ( .A(n3082), .B(n3077), .C(n3078), .D(n3083), .Y(n_1609) );
    zoai22d U1234 ( .A(n3084), .B(n3077), .C(n3078), .D(n3085), .Y(n_1611) );
    zoai22d U1235 ( .A(n3087), .B(n3077), .C(n3078), .D(n3088), .Y(n_1615) );
    zoai22d U1236 ( .A(n3089), .B(n3090), .C(n3091), .D(n3092), .Y(n_1236) );
    zoai22d U1237 ( .A(n3093), .B(n3090), .C(n3091), .D(n3094), .Y(n_1238) );
    zoai22d U1238 ( .A(n3095), .B(n3090), .C(n3091), .D(n3096), .Y(n_1240) );
    zoai22d U1239 ( .A(n3097), .B(n3090), .C(n3091), .D(n3098), .Y(n_1242) );
    zao222b U1240 ( .A(n3099), .B(AD3I), .C(n2983), .D(ENUSB4), .E(HCSPARAMS_3
        ), .F(n3100), .Y(n_1244) );
    zao222b U1241 ( .A(n3099), .B(AD2I), .C(n2983), .D(n2980), .E(HCSPARAMS_2), 
        .F(n3100), .Y(n_1246) );
    zao222b U1242 ( .A(n3099), .B(AD1I), .C(n2983), .D(n2981), .E(HCSPARAMS_1), 
        .F(n3100), .Y(n_1248) );
    zoai22d U1243 ( .A(n3101), .B(n3090), .C(n3091), .D(n3102), .Y(n_1250) );
    zoai22d U1244 ( .A(n3103), .B(n3104), .C(n3105), .D(n3106), .Y(
        FRLSTSIZE1579_0) );
    zoai22d U1245 ( .A(n3103), .B(n3107), .C(n3108), .D(n3109), .Y(
        FRLSTSIZE1579_1) );
    zor5b U1246 ( .A(n3110), .B(n3111), .C(n3112), .D(n3113), .E(n3114), .Y(
        REGDOUT2[0]) );
    zor4b U1247 ( .A(n3115), .B(n3116), .C(n3117), .D(n3118), .Y(REGDOUT2[1])
         );
    zor4b U1248 ( .A(n3119), .B(n3120), .C(n3121), .D(n3122), .Y(REGDOUT2[2])
         );
    zor4b U1249 ( .A(n3123), .B(n3124), .C(n3125), .D(n3126), .Y(REGDOUT2[3])
         );
    zor6b U1250 ( .A(n3127), .B(n3128), .C(n3129), .D(n3130), .E(n3131), .F(
        n3132), .Y(REGDOUT2[4]) );
    zor4b U1251 ( .A(n3133), .B(n3134), .C(n3135), .D(n3136), .Y(REGDOUT2[5])
         );
    zor6b U1252 ( .A(n3137), .B(n3138), .C(n3139), .D(n3140), .E(n3141), .F(
        n3142), .Y(REGDOUT2[6]) );
    zor6b U1253 ( .A(n3143), .B(n3144), .C(n3145), .D(n3146), .E(n3147), .F(
        n3148), .Y(REGDOUT2[7]) );
    zor4b U1254 ( .A(n3169), .B(n3170), .C(n3171), .D(n3172), .Y(REGDOUT2[12])
         );
    zor4b U1255 ( .A(n3173), .B(n3174), .C(n3175), .D(n3176), .Y(REGDOUT2[13])
         );
    zor6b U1256 ( .A(n3177), .B(n3178), .C(n3179), .D(n3180), .E(n3181), .F(
        n3182), .Y(REGDOUT2[14]) );
    zor6b U1257 ( .A(n3183), .B(n3184), .C(n3185), .D(n3186), .E(n3187), .F(
        n3188), .Y(REGDOUT2[15]) );
    zor6b U1258 ( .A(n3209), .B(n3210), .C(n3211), .D(n3212), .E(n3213), .F(
        n3214), .Y(REGDOUT2[20]) );
    zor3b U1259 ( .A(n3230), .B(n3231), .C(n3232), .Y(REGDOUT2[24]) );
    zor3b U1260 ( .A(n3233), .B(n3234), .C(n3235), .Y(REGDOUT2[25]) );
    zor3b U1261 ( .A(n3236), .B(n3237), .C(n3238), .Y(REGDOUT2[26]) );
    zor3b U1262 ( .A(n3239), .B(n3240), .C(n3241), .Y(REGDOUT2[27]) );
    zor3b U1263 ( .A(n3242), .B(n3243), .C(n3244), .Y(REGDOUT2[28]) );
    zor3b U1264 ( .A(n3245), .B(n3246), .C(n3247), .Y(REGDOUT2[29]) );
    zor3b U1265 ( .A(n3248), .B(n3249), .C(n3250), .Y(REGDOUT2[30]) );
    zor3b U1266 ( .A(n3251), .B(n3252), .C(n3253), .Y(REGDOUT2[31]) );
    zoa21d U1267 ( .A(ENUSB2), .B(n3255), .C(n3256), .Y(n3254) );
    zoa21d U1268 ( .A(n3257), .B(n3258), .C(USBLEGCTLSTS[29]), .Y(n3038) );
    zoa21d U1269 ( .A(n3109), .B(n3259), .C(USBLEGCTLSTS[19]), .Y(n3039) );
    zoa21d U1270 ( .A(n3106), .B(n3259), .C(USBLEGCTLSTS[18]), .Y(n3040) );
    zoa21d U1271 ( .A(n3097), .B(n3259), .C(USBLEGCTLSTS[20]), .Y(n3041) );
    zoa21d U1272 ( .A(n3260), .B(n3258), .C(USBLEGCTLSTS[31]), .Y(n3042) );
    zoa21d U1273 ( .A(n3261), .B(n3259), .C(ERRINT), .Y(n3043) );
    zoa21d U1274 ( .A(n3095), .B(n3259), .C(INTASYNC), .Y(n3034) );
    zoa21d U1275 ( .A(n3101), .B(n3259), .C(USBINT), .Y(n3036) );
    zoa21d U1276 ( .A(n3262), .B(n3258), .C(USBLEGCTLSTS[30]), .Y(n3035) );
    zoa21d U1277 ( .A(AD2I), .B(n3264), .C(n3107), .Y(n3108) );
    zoa21d U1278 ( .A(AD3I), .B(n3264), .C(n3104), .Y(n3105) );
    zor3b U1279 ( .A(PA4I), .B(PA7I), .C(PA6I), .Y(n3269) );
    zor4b U1280 ( .A(n3324), .B(n3325), .C(n3326), .D(n3327), .Y(n3323) );
    zor2d U1281 ( .A(n3080), .B(n3323), .Y(n3078) );
    zor3b U1282 ( .A(n3275), .B(n3321), .C(n3296), .Y(n3077) );
    zor3b U1283 ( .A(n3270), .B(n3275), .C(n3332), .Y(n3090) );
    zor3b U1284 ( .A(PA6I), .B(PA5I), .C(n3336), .Y(n3338) );
    zor4b U1285 ( .A(CBE3I_), .B(CBE0I_), .C(CBE1I_), .D(n3284), .Y(n3339) );
    zor3b U1286 ( .A(n3269), .B(n3340), .C(n3339), .Y(n3341) );
    zor4b U1287 ( .A(PA4I), .B(PA6I), .C(n3367), .D(n3340), .Y(n3368) );
    zor4b U1288 ( .A(n3340), .B(n3367), .C(PA6I), .D(n3335), .Y(n3374) );
    zor3b U1289 ( .A(n3378), .B(n3340), .C(n3336), .Y(n3379) );
    zor4b U1290 ( .A(PA4I), .B(PA7I), .C(n3378), .D(n3340), .Y(n3381) );
    zor3b U1291 ( .A(PA5I), .B(n3378), .C(n3336), .Y(n3386) );
    zor3b U1292 ( .A(n3340), .B(n3295), .C(n3269), .Y(n3390) );
    zor3b U1293 ( .A(n3340), .B(n3320), .C(n3269), .Y(n3396) );
    zao333b U1294 ( .A(USBLEGCTLSTS[0]), .B(n3358), .C(USBINT_S), .D(
        USBLEGCTLSTS[14]), .E(n3365), .F(PCI_RPCMD), .G(USBLEGCTLSTS[13]), .H(
        n3342), .I(SMIOSOWNCHG_NXT), .Y(n3032) );
    zao222b U1295 ( .A(PORTCHG_EN), .B(USBLEGCTLSTS[18]), .C(HSERR_EN), .D(
        USBLEGCTLSTS[20]), .E(ROLLOVER_EN), .F(USBLEGCTLSTS[19]), .Y(n3064) );
    zind2d U1296 ( .A(INTR_DIS), .B(PWR_STATE_D0), .Y(n3071) );
    zor3b U1297 ( .A(TABORTR), .B(RUN_C), .C(HCRESET), .Y(n3446) );
    zao222b U1298 ( .A(DBGPORT_SC[7]), .B(n2996), .C(DBGPORT_PID[7]), .D(n3069
        ), .E(DBGPORT_BUF2[7]), .F(n3448), .Y(n3148) );
    zao222b U1299 ( .A(PORTSC2[7]), .B(n3510), .C(PORTSC4[7]), .D(n3063), .E(
        PORTSC3[7]), .F(n3009), .Y(n3145) );
    zao222b U1300 ( .A(DBGPORT_SC[6]), .B(n2995), .C(DBGPORT_PID[6]), .D(n2990
        ), .E(DBGPORT_BUF2[6]), .F(n3448), .Y(n3142) );
    zao222b U1301 ( .A(PORTSC2[6]), .B(n3510), .C(PORTSC4[6]), .D(n3063), .E(
        PORTSC3[6]), .F(n3507), .Y(n3139) );
    zao222b U1302 ( .A(DBGPORT_SC[5]), .B(n2995), .C(DBGPORT_PID[5]), .D(n2989
        ), .E(DBGPORT_BUF2[5]), .F(n3514), .Y(n3453) );
    zao222b U1303 ( .A(PORTSC6[5]), .B(n3008), .C(PORTSC8[5]), .D(n3067), .E(
        PORTSC7[5]), .F(n3050), .Y(n3133) );
    zor5b U1304 ( .A(n3454), .B(n3455), .C(n3456), .D(n3457), .E(n3453), .Y(
        n3136) );
    zao222b U1305 ( .A(FRNUM_SYNC_5), .B(n2979), .C(ASYNCLISTADDR[5]), .D(
        n3449), .E(PORTSC3[5]), .F(n3062), .Y(n3456) );
    zao222b U1306 ( .A(n3452), .B(ASYNC_EN), .C(n3459), .D(INTASYNC), .E(
        HCSPARAMS_5), .F(n3451), .Y(n3454) );
    zao222b U1307 ( .A(DBGPORT_PID[4]), .B(n2990), .C(DBGPORT_ADDR[4]), .D(
        n3056), .E(DBGPORT_BUF2[4]), .F(n3448), .Y(n3132) );
    zao211b U1308 ( .A(DBGPORT_BUF1[4]), .B(n3447), .C(n3460), .D(n3461), .Y(
        n3131) );
    zao222b U1309 ( .A(PORTSC5[4]), .B(n3005), .C(PORTSC6[4]), .D(n3512), .E(
        DBGPORT_SC[4]), .F(n3505), .Y(n3462) );
    zao211b U1310 ( .A(PORTSC8[4]), .B(n2992), .C(n3263), .D(n3462), .Y(n3461)
         );
    zao222b U1311 ( .A(PORTSC2[4]), .B(n3510), .C(PORTSC4[4]), .D(n3063), .E(
        PORTSC3[4]), .F(n3009), .Y(n3129) );
    zao222b U1312 ( .A(n3452), .B(PERIOD_EN), .C(n3459), .D(USBLEGCTLSTS[20]), 
        .E(HCSPARAMS_4), .F(n3451), .Y(n3127) );
    zao222b U1313 ( .A(DBGPORT_PID[31]), .B(n2989), .C(DBGPORT_ADDR[31]), .D(
        n3506), .E(DBGPORT_BUF1[31]), .F(n3513), .Y(n3463) );
    zao211b U1314 ( .A(DBGPORT_BUF2[31]), .B(n3448), .C(n3464), .D(n3463), .Y(
        n3253) );
    zao222b U1315 ( .A(DBGPORT_PID[30]), .B(n2990), .C(DBGPORT_ADDR[30]), .D(
        n3003), .E(DBGPORT_BUF1[30]), .F(n3447), .Y(n3466) );
    zao211b U1316 ( .A(DBGPORT_BUF2[30]), .B(n3514), .C(n3467), .D(n3466), .Y(
        n3250) );
    zao222b U1317 ( .A(DBGPORT_SC[3]), .B(n2996), .C(DBGPORT_PID[3]), .D(n2989
        ), .E(DBGPORT_BUF2[3]), .F(n3514), .Y(n3468) );
    zao222b U1318 ( .A(PORTSC6[3]), .B(n3059), .C(PORTSC8[3]), .D(n2992), .E(
        PORTSC7[3]), .F(n3050), .Y(n3123) );
    zor4b U1319 ( .A(n3469), .B(n3470), .C(n3471), .D(n3468), .Y(n3126) );
    zao222b U1320 ( .A(FRLSTSIZE[1]), .B(n3452), .C(FRNUM_SYNC_3), .D(n2979), 
        .E(PORTSC3[3]), .F(n3062), .Y(n3469) );
    zao222b U1321 ( .A(DBGPORT_PID[29]), .B(n2990), .C(DBGPORT_ADDR[29]), .D(
        n3506), .E(DBGPORT_BUF1[29]), .F(n3513), .Y(n3472) );
    zao211b U1322 ( .A(DBGPORT_BUF2[29]), .B(n3448), .C(n3473), .D(n3472), .Y(
        n3247) );
    zao222b U1323 ( .A(DBGPORT_PID[28]), .B(n2989), .C(DBGPORT_ADDR[28]), .D(
        n3056), .E(DBGPORT_BUF1[28]), .F(n3447), .Y(n3474) );
    zao211b U1324 ( .A(DBGPORT_BUF2[28]), .B(n3514), .C(n3475), .D(n3474), .Y(
        n3244) );
    zao222b U1325 ( .A(DBGPORT_PID[27]), .B(n3069), .C(DBGPORT_ADDR[27]), .D(
        n3506), .E(DBGPORT_BUF1[27]), .F(n3513), .Y(n3476) );
    zao211b U1326 ( .A(DBGPORT_BUF2[27]), .B(n3448), .C(n3477), .D(n3476), .Y(
        n3241) );
    zao222b U1327 ( .A(DBGPORT_PID[26]), .B(n3069), .C(DBGPORT_ADDR[26]), .D(
        n3056), .E(DBGPORT_BUF1[26]), .F(n3447), .Y(n3478) );
    zao211b U1328 ( .A(DBGPORT_BUF2[26]), .B(n3514), .C(n3479), .D(n3478), .Y(
        n3238) );
    zao222b U1329 ( .A(DBGPORT_PID[25]), .B(n2989), .C(DBGPORT_ADDR[25]), .D(
        n3506), .E(DBGPORT_BUF1[25]), .F(n3513), .Y(n3480) );
    zao211b U1330 ( .A(DBGPORT_BUF2[25]), .B(n3448), .C(n3481), .D(n3480), .Y(
        n3235) );
    zao222b U1331 ( .A(DBGPORT_PID[24]), .B(n3069), .C(DBGPORT_ADDR[24]), .D(
        n3056), .E(DBGPORT_BUF1[24]), .F(n3447), .Y(n3482) );
    zao211b U1332 ( .A(DBGPORT_BUF2[24]), .B(n3514), .C(n3483), .D(n3482), .Y(
        n3232) );
    zao222b U1333 ( .A(DBGPORT_SC[20]), .B(n3505), .C(DBGPORT_PID[20]), .D(
        n2989), .E(DBGPORT_BUF2[20]), .F(n3448), .Y(n3214) );
    zao222b U1334 ( .A(PORTSC2[20]), .B(n3510), .C(PORTSC4[20]), .D(n2999), 
        .E(PORTSC3[20]), .F(n3009), .Y(n3209) );
    zao222b U1335 ( .A(DBGPORT_SC[2]), .B(n2996), .C(DBGPORT_PID[2]), .D(n2990
        ), .E(DBGPORT_BUF2[2]), .F(n3514), .Y(n3484) );
    zao222b U1336 ( .A(PORTSC6[2]), .B(n3008), .C(PORTSC8[2]), .D(n2993), .E(
        PORTSC7[2]), .F(n3010), .Y(n3119) );
    zor4b U1337 ( .A(n3485), .B(n3486), .C(n3487), .D(n3484), .Y(n3122) );
    zao222b U1338 ( .A(FRLSTSIZE[0]), .B(n3452), .C(FRNUM_SYNC_2), .D(n2979), 
        .E(PORTSC3[2]), .F(n3062), .Y(n3485) );
    zao222b U1339 ( .A(DBGPORT_SC[15]), .B(n2995), .C(DBGPORT_PID[15]), .D(
        n2990), .E(DBGPORT_BUF2[15]), .F(n3448), .Y(n3188) );
    zao222b U1340 ( .A(PORTSC2[15]), .B(n3007), .C(PORTSC4[15]), .D(n2998), 
        .E(PORTSC3[15]), .F(n3009), .Y(n3185) );
    zao222b U1341 ( .A(DBGPORT_SC[14]), .B(n3505), .C(DBGPORT_PID[14]), .D(
        n3069), .E(DBGPORT_BUF2[14]), .F(n3514), .Y(n3182) );
    zao222b U1342 ( .A(PORTSC2[14]), .B(n3007), .C(PORTSC4[14]), .D(n2998), 
        .E(PORTSC3[14]), .F(n3507), .Y(n3179) );
    zao222b U1343 ( .A(DBGPORT_SC[13]), .B(n2995), .C(DBGPORT_PID[13]), .D(
        n3069), .E(DBGPORT_BUF2[13]), .F(n3448), .Y(n3488) );
    zao222b U1344 ( .A(PORTSC6[13]), .B(n3008), .C(PORTSC8[13]), .D(n2993), 
        .E(PORTSC7[13]), .F(n3010), .Y(n3173) );
    zor4b U1345 ( .A(n3489), .B(n3490), .C(n3491), .D(n3488), .Y(n3176) );
    zao222b U1346 ( .A(FRNUM_SYNC_13), .B(n2979), .C(ASYNCLISTADDR[13]), .D(
        n3449), .E(PORTSC3[13]), .F(n3062), .Y(n3489) );
    zao222b U1347 ( .A(DBGPORT_SC[12]), .B(n2995), .C(DBGPORT_PID[12]), .D(
        n3069), .E(DBGPORT_BUF2[12]), .F(n3514), .Y(n3492) );
    zao222b U1348 ( .A(PORTSC6[12]), .B(n3059), .C(PORTSC8[12]), .D(n2992), 
        .E(PORTSC7[12]), .F(n3010), .Y(n3169) );
    zor4b U1349 ( .A(n3493), .B(n3494), .C(n3495), .D(n3492), .Y(n3172) );
    zao222b U1350 ( .A(FRNUM_SYNC_12), .B(n2979), .C(ASYNCLISTADDR[12]), .D(
        n3449), .E(PORTSC3[12]), .F(n3062), .Y(n3493) );
    zao222b U1351 ( .A(DBGPORT_SC[1]), .B(n2995), .C(DBGPORT_PID[1]), .D(n2989
        ), .E(DBGPORT_BUF2[1]), .F(n3448), .Y(n3496) );
    zao222b U1352 ( .A(PORTSC6[1]), .B(n3059), .C(PORTSC8[1]), .D(n3067), .E(
        PORTSC7[1]), .F(n3010), .Y(n3115) );
    zor4b U1353 ( .A(n3497), .B(n3498), .C(n3499), .D(n3496), .Y(n3118) );
    zao222b U1354 ( .A(HCSPARAMS_1), .B(n3451), .C(FRNUM_SYNC_1), .D(n2979), 
        .E(PORTSC3[1]), .F(n3062), .Y(n3499) );
    zao222b U1355 ( .A(DBGPORT_PID[0]), .B(n3069), .C(DBGPORT_ADDR[0]), .D(
        n3506), .E(DBGPORT_BUF2[0]), .F(n3514), .Y(n3501) );
    zao222b U1356 ( .A(PORTSC5[0]), .B(n3511), .C(PORTSC6[0]), .D(n3512), .E(
        DBGPORT_SC[0]), .F(n2996), .Y(n3503) );
    zor4b U1357 ( .A(n3503), .B(n3502), .C(n3500), .D(n3501), .Y(n3114) );
    zao222b U1358 ( .A(PORTSC2[0]), .B(n3007), .C(PORTSC4[0]), .D(n2998), .E(
        PORTSC3[0]), .F(n3507), .Y(n3112) );
    zao222b U1359 ( .A(RUN), .B(n3452), .C(n3459), .D(USBINT), .E(HCSPARAMS_0), 
        .F(n3451), .Y(n3110) );
    zan2d S_4 ( .A(HRST_), .B(n_12), .Y(n_13) );
    zan2d S_6 ( .A(n_13), .B(n_14), .Y(n_15) );
    zor2d S_7 ( .A(n_15), .B(ATPG_ENI), .Y(n3526) );
    zbfb U1360 ( .A(HCRESET), .Y(n3517) );
    zbfb U1361 ( .A(USMIACT_T), .Y(n3518) );
    zbfb U1362 ( .A(LIGHTRST), .Y(n3519) );
    zbfb U1363 ( .A(USMIO_T), .Y(n3520) );
    zbfb U1364 ( .A(LIGHTRST_T), .Y(n3521) );
    zbfb U1365 ( .A(HCRESET_T), .Y(n3522) );
    zbfp U1366 ( .A(n3526), .Y(CMDRST_) );
    zbfp U1367 ( .A(n3526), .Y(n3524) );
    zbfp U1368 ( .A(n3526), .Y(n3525) );
endmodule


module HS_PCICFG ( CFGD31, CFGD30, CFGD29, CFGD28, CFGD27, CFGD26, CFGD25, 
    CFGD24, CFGD23, CFGD22, CFGD21, CFGD20, CFGD19, CFGD18, CFGD17, CFGD16, 
    CFGD15, CFGD14, CFGD13, CFGD12, CFGD11, CFGD10, CFGD9, CFGD8, CFGD7, CFGD6, 
    CFGD5, CFGD4, CFGD3, CFGD2, CFGD1, CFGD0, IOBA31, IOBA30, IOBA29, IOBA28, 
    IOBA27, IOBA26, IOBA25, IOBA24, IOBA23, IOBA22, IOBA21, IOBA20, IOBA19, 
    IOBA18, IOBA17, IOBA16, IOBA15, IOBA14, IOBA13, IOBA12, IOBA11, IOBA10, 
    IOBA9, IOBA8, CACHLN7, CACHLN6, CACHLN5, CACHLN4, CACHLN3, CACHLN2, 
    CACHLN1, CACHLN0, DEVS0, INTR_DIS, FB2BKEN, SERREN, RSTEP, RPTYERR, MWRMEN, 
    BMASTREN, MMSPACE, IOSPACE, UIRQSEL3, UIRQSEL2, UIRQSEL1, UIRQSEL0, 
    PCI1WAIT, FCFG, PM_EN, HCISPEC_, REDUCE, PAROPT, BABOPT, CAHCFG_, TRAP_OPT, 
    VIAPSS, DBGIRQ, TESTCNT, ENOCPY, DISEOP, DISPRST, DISSTUFF, RxDataOut_A, 
    SquelchOut_A, DisconnectOut_A, TERM_ON_A, RxDataOut_B, SquelchOut_B, 
    DisconnectOut_B, TERM_ON_B, RxDataOut_C, SquelchOut_C, DisconnectOut_C, 
    TERM_ON_C, RxDataOut_D, SquelchOut_D, DisconnectOut_D, TERM_ON_D, 
    RxDataOut_E, SquelchOut_E, DisconnectOut_E, TERM_ON_E, RxDataOut_F, 
    SquelchOut_F, DisconnectOut_F, TERM_ON_F, RxDataOut_G, SquelchOut_G, 
    DisconnectOut_G, TERM_ON_G, RxDataOut_H, SquelchOut_H, DisconnectOut_H, 
    TERM_ON_H, AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I, AD23I, 
    AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, AD14I, AD13I, 
    AD12I, AD11I, AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, 
    AD0I, PA7I, PA6I, PA5I, PA4I, PA3I, PA2I, CBE3I_, CBE2I_, CBE1I_, CBE0I_, 
    CFGW, FLADJ5, FLADJ4, FLADJ3, FLADJ2, FLADJ1, FLADJ0, PORTWAKECAP8, 
    PORTWAKECAP7, PORTWAKECAP6, PORTWAKECAP5, PORTWAKECAP4, PORTWAKECAP3, 
    PORTWAKECAP2, PORTWAKECAP1, PORTWAKECAP0, PME_EN, PME_STS, PWR_STATE1, 
    PWR_STATE0, E_PME_EN, EN_DBG_PORT, R61G, R62G, R63G, R84G, R85G, PCI_R6AG, 
    PCI_R6BG, PCI_R6CG, PCI_R6DG, PCI_R6FG, PCI_RBAR, PCI_RPCMD, REVID7, 
    REVID6, REVID5, REVID4, REVID3, REVID2, REVID1, REVID0, MAXLAT7, MAXLAT6, 
    MAXLAT5, MAXLAT4, MAXLAT3, MAXLAT2, MAXLAT1, MAXLAT0, MINGNT7, MINGNT6, 
    MINGNT5, MINGNT4, MINGNT3, MINGNT2, MINGNT1, MINGNT0, UIRQACT, SERRS, 
    MABORTS, TABORTR, OCUPY_SEL, DISTXDLY, DISPFUNDRN, ENTXDLY_1, ENTXDLY_2, 
    ENTXDLY_3, SELEOF, DISTXDLY2, DISFFCRC0, DISFFCRC1, DISPFIFO, DISPFIFO2, 
    DISRXZERO, ENBMUSMRST, FUNCSEL, DISPSTUFF, SLQUEUEADDR, SWDBG, SLAVEMODE, 
    SLAVE_ACT, SL_ERROFFSET, CRCERR, PIDERR, SL_DATA_PIDERR, SL_ET_ERR, 
    SL_SE_ERR, SL_ACK_ERR, SL_PCIERR, SLAVE_ERR, BIST_RUN, BIST_RUN_C, 
    BIST_ERR_S, DIS_BURST, TMOUT_PARM, ENISOHANDCHK, DISCHKEOPERR, HCHALT, 
    CMDRST_, CP0, CP1, SOF_DISCONN_CHK, CTRL_A, CTRL_B, CTRL_C, CTRL_D, CTRL_E, 
    CTRL_F, CTRL_G, CTRL_H, tst_buferr, loopback, tstmod, rx_block_dis, 
    FastLock, LockSpd, TrkSpd, RxDataDly, FastStart, autochk, sync_fast, 
    sync_jend, SQSET, RDOUT_Enb, LBack_Enb, FAST_RST, TMODE, BypassDiv4, 
    UTM_CHKERR, TEST_EYE_EN, FORCE_CRCERR, DIS_NARROW_SOF, SetPowner_Dis, 
    PdPHY_Dis, HsEnFB_Dis, DIS_TERM_ON_A, DIS_TERM_ON_B, DIS_TERM_ON_C, 
    DIS_TERM_ON_D, DIS_TERM_ON_E, DIS_TERM_ON_F, DIS_TERM_ON_G, DIS_TERM_ON_H, 
    USBLEGCTLSTS, USBLEGSUP, SUBIDWE, DISPDRCV, CLKOFF_EN, TXTMOUT_EN, 
    TXDELAY_EN, TXDELAY_PARM, TURN_PARM, ENUSB1, ENUSB2, ENUSB3, ENUSB4, 
    DIS_SOF_RUN, SLEEPTIME_SEL, BIST_PATTERN, SRAM_WR, SRAM_RUN, SRAM_ADDR, 
    SRAM_SEL, SRAM_RDATA1, SRAM_RDATA2, SRAM_RDATA3, SRAM_RDATA4, EN_CHKTOGCRC, 
    EN_UTM_RESET, EN_REF_RVLD, EN_UTM_SPDUP, PCICLK, PCICLK_FREE, HRST_ );
output [1:0] OCUPY_SEL;
input  [2:0] FUNCSEL;
output [3:0] CTRL_H;
output [1:0] LockSpd;
output [31:0] SLQUEUEADDR;
input  [7:0] SL_ERROFFSET;
output [3:0] CTRL_A;
output [3:0] CTRL_F;
output [1:0] SQSET;
input  [31:0] SRAM_RDATA2;
output [3:0] CTRL_G;
output [3:0] TURN_PARM;
output [31:0] BIST_PATTERN;
output [8:0] SRAM_ADDR;
input  [31:0] SRAM_RDATA3;
output [3:0] CTRL_B;
output [1:0] TrkSpd;
input  [31:0] USBLEGSUP;
input  [31:0] SRAM_RDATA4;
output [3:0] CTRL_D;
output [3:0] CTRL_E;
output [2:0] RxDataDly;
output [7:0] TXDELAY_PARM;
input  [31:0] SRAM_RDATA1;
input  [31:0] USBLEGCTLSTS;
output [7:0] TMOUT_PARM;
output [3:0] CTRL_C;
output [1:0] SRAM_SEL;
input  RxDataOut_A, SquelchOut_A, DisconnectOut_A, TERM_ON_A, RxDataOut_B, 
    SquelchOut_B, DisconnectOut_B, TERM_ON_B, RxDataOut_C, SquelchOut_C, 
    DisconnectOut_C, TERM_ON_C, RxDataOut_D, SquelchOut_D, DisconnectOut_D, 
    TERM_ON_D, RxDataOut_E, SquelchOut_E, DisconnectOut_E, TERM_ON_E, 
    RxDataOut_F, SquelchOut_F, DisconnectOut_F, TERM_ON_F, RxDataOut_G, 
    SquelchOut_G, DisconnectOut_G, TERM_ON_G, RxDataOut_H, SquelchOut_H, 
    DisconnectOut_H, TERM_ON_H, AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, 
    AD25I, AD24I, AD23I, AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I, 
    AD15I, AD14I, AD13I, AD12I, AD11I, AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, 
    AD4I, AD3I, AD2I, AD1I, AD0I, PA7I, PA6I, PA5I, PA4I, PA3I, PA2I, CBE3I_, 
    CBE2I_, CBE1I_, CBE0I_, CFGW, FLADJ5, FLADJ4, FLADJ3, FLADJ2, FLADJ1, 
    FLADJ0, PORTWAKECAP8, PORTWAKECAP7, PORTWAKECAP6, PORTWAKECAP5, 
    PORTWAKECAP4, PORTWAKECAP3, PORTWAKECAP2, PORTWAKECAP1, PORTWAKECAP0, 
    PME_EN, PME_STS, PWR_STATE1, PWR_STATE0, E_PME_EN, REVID7, REVID6, REVID5, 
    REVID4, REVID3, REVID2, REVID1, REVID0, MAXLAT7, MAXLAT6, MAXLAT5, MAXLAT4, 
    MAXLAT3, MAXLAT2, MAXLAT1, MAXLAT0, MINGNT7, MINGNT6, MINGNT5, MINGNT4, 
    MINGNT3, MINGNT2, MINGNT1, MINGNT0, UIRQACT, SERRS, MABORTS, TABORTR, 
    SLAVE_ACT, CRCERR, PIDERR, SL_DATA_PIDERR, SL_ET_ERR, SL_SE_ERR, 
    SL_ACK_ERR, SL_PCIERR, SLAVE_ERR, BIST_RUN_C, BIST_ERR_S, HCHALT, CMDRST_, 
    UTM_CHKERR, ENUSB1, ENUSB2, ENUSB3, ENUSB4, PCICLK, PCICLK_FREE, HRST_;
output CFGD31, CFGD30, CFGD29, CFGD28, CFGD27, CFGD26, CFGD25, CFGD24, CFGD23, 
    CFGD22, CFGD21, CFGD20, CFGD19, CFGD18, CFGD17, CFGD16, CFGD15, CFGD14, 
    CFGD13, CFGD12, CFGD11, CFGD10, CFGD9, CFGD8, CFGD7, CFGD6, CFGD5, CFGD4, 
    CFGD3, CFGD2, CFGD1, CFGD0, IOBA31, IOBA30, IOBA29, IOBA28, IOBA27, IOBA26, 
    IOBA25, IOBA24, IOBA23, IOBA22, IOBA21, IOBA20, IOBA19, IOBA18, IOBA17, 
    IOBA16, IOBA15, IOBA14, IOBA13, IOBA12, IOBA11, IOBA10, IOBA9, IOBA8, 
    CACHLN7, CACHLN6, CACHLN5, CACHLN4, CACHLN3, CACHLN2, CACHLN1, CACHLN0, 
    DEVS0, INTR_DIS, FB2BKEN, SERREN, RSTEP, RPTYERR, MWRMEN, BMASTREN, 
    MMSPACE, IOSPACE, UIRQSEL3, UIRQSEL2, UIRQSEL1, UIRQSEL0, PCI1WAIT, FCFG, 
    PM_EN, HCISPEC_, REDUCE, PAROPT, BABOPT, CAHCFG_, TRAP_OPT, VIAPSS, DBGIRQ, 
    TESTCNT, ENOCPY, DISEOP, DISPRST, DISSTUFF, EN_DBG_PORT, R61G, R62G, R63G, 
    R84G, R85G, PCI_R6AG, PCI_R6BG, PCI_R6CG, PCI_R6DG, PCI_R6FG, PCI_RBAR, 
    PCI_RPCMD, DISTXDLY, DISPFUNDRN, ENTXDLY_1, ENTXDLY_2, ENTXDLY_3, SELEOF, 
    DISTXDLY2, DISFFCRC0, DISFFCRC1, DISPFIFO, DISPFIFO2, DISRXZERO, 
    ENBMUSMRST, DISPSTUFF, SWDBG, SLAVEMODE, BIST_RUN, DIS_BURST, ENISOHANDCHK, 
    DISCHKEOPERR, CP0, CP1, SOF_DISCONN_CHK, tst_buferr, loopback, tstmod, 
    rx_block_dis, FastLock, FastStart, autochk, sync_fast, sync_jend, 
    RDOUT_Enb, LBack_Enb, FAST_RST, TMODE, BypassDiv4, TEST_EYE_EN, 
    FORCE_CRCERR, DIS_NARROW_SOF, SetPowner_Dis, PdPHY_Dis, HsEnFB_Dis, 
    DIS_TERM_ON_A, DIS_TERM_ON_B, DIS_TERM_ON_C, DIS_TERM_ON_D, DIS_TERM_ON_E, 
    DIS_TERM_ON_F, DIS_TERM_ON_G, DIS_TERM_ON_H, SUBIDWE, DISPDRCV, CLKOFF_EN, 
    TXTMOUT_EN, TXDELAY_EN, DIS_SOF_RUN, SLEEPTIME_SEL, SRAM_WR, SRAM_RUN, 
    EN_CHKTOGCRC, EN_UTM_RESET, EN_REF_RVLD, EN_UTM_SPDUP;
    wire RxData_B, IOBA292419, n_10876, n_5138, DEBUGB3287_5, PHYOPT13477_5, 
        DEBUGD3363_0, TMABORTS, PHYMON_EN_F4392, SUBSID0_4, MMSPACE2040, 
        n_8054, SUBVID12860_1, TERMON_C, Squelch_H, PHYOPT43591_1, 
        LAT_TM2299_7, IOBA162538, SPAREO6, DEBUG02974_0, DEBUG23050_5, 
        INTLN2337_1, REVID_BACK_2, SUBSID12936_2, CACHLN02164, DEBUGF_3, 
        Disconnect_E, SRAM_RDATA_SEL_2, SUBSID1_4, RxDataDly3781_2, 
        PHYOPT33553_6, IOBA112705, DEBUGA3249_0, BIST_ERROR4199, BMASTREN2046, 
        n_5660, TMOUT_PARM4236_2, n_10888, n_6198, PHYOPTGH3667_0, 
        Disconnect_G5019, SRAM_RDATA_SEL_11, SRAM_RUN_T, IOBA102699, 
        TERMON_H5098, SRAM_RDATA_SEL_24, SRAM_ADDR_IN_7, DEBUG83126_2, n_9566, 
        BACK_EN, Squelch_A, n_5672, DEBUG33088_6, DEBUGC3325_3, INTLN_2, 
        PHYMON_EN_C, SRAM_SEL5343_0, DEBUGF3439_4, IOBA312431, DEBUG13012_5, 
        DEBUGD_6, n_8046, n_2808, DEBUGE3401_4, SUBVID02822_5, RxData_D4776, 
        SUBSID02898_3, REVID_BACK5677_7, INTR_DIS2113, PHYOPTEF3629_2, 
        Disconnect_D4764, MWRMEN2052, n_10220, SRAM_RDATA_SEL_18, 
        PHYOPT23515_4, CACHLN32182, IOBA242389, n_6196, SUBSID02898_4, 
        SUBVID02822_2, DEBUGE3401_3, PHYOPT23515_3, SUBVID0_0, PHYOPTEF3629_5, 
        CACHLN42188, REVID_BACK5677_0, DEBUG13012_2, DEBUGF3439_3, PHYMON_EN_D, 
        SPAREO0_, n_10886, DEBUGC3325_4, DEBUG33088_1, Squelch_F, DEBUGE_1, 
        SPAREO8, TERMON_C4673, TrkSpd3743_1, n_6730, SRAM_ADDR_IN_0, 
        SRAM_RDATA_SEL_23, n_10878, n_5136, SUBVID1_0, n_11542, DEBUG83126_5, 
        Squelch_D4770, PHYOPTGH3667_7, n_11550, n_6722, SRAM_RDATA_SEL_31, 
        TERMON_F4928, SRAM_RDATA_SEL_16, SRAM_RDATA_SEL_5, Disconnect_B, 
        DEBUGB3287_2, SUBSID12936_5, n_8048, TMOUT_PARM4236_5, n_2806, 
        DEBUGA3249_7, PHYOPT33553_1, PHYOPT43591_6, CACHLN62200, TERMON_D, 
        SUBVID12860_6, SUBSID0_3, REVID_BACK_5, INTLN2337_6, DEBUG23050_2, 
        DEBUG02974_7, SPAREO1, LAT_TM2299_0, IOBA232580, RxData_E, n_9568, 
        SRAM_RUN5389, DEBUGD3363_7, PHYOPT13477_2, Squelch_F4940, 
        SRAM_RDATA_SEL_22, SRAM_ADDR_IN_1, INTLN_4, CACHLN22176, DEBUG83126_4, 
        IOBA132717, n_9560, IOBA182550, DEBUGC3325_5, DEBUG33088_0, Squelch_G, 
        SPAREO9, TrkSpd3743_0, DEBUG13012_3, DEBUGF3439_2, n_5142, PHYMON_EN_E, 
        TERMON_D4758, n_11536, PHYMON_EN_D4380, n_8040, SUBSID02898_5, 
        FB2BKENR, SUBVID02822_3, DEBUGE3401_2, FBCYC, PHYOPT23515_2, SUBVID0_1, 
        n_10226, REVID_BACK5677_1, PHYOPTEF3629_4, FORCE_CRCERR4311, 
        SRAM_ADDR_IN_8, SWDBG4088, RxData_D, RxData_G5031, DEBUGB3287_3, 
        DEBUGD3363_6, PHYOPT13477_3, RxData_C4691, PHYOPT43591_7, TERMON_E, 
        IOBA282413, n_8052, SUBVID12860_7, SUBSID0_2, INTLN2337_7, 
        REVID_BACK_4, DEBUG23050_3, DEBUG02974_6, SPAREO0, LAT_TM2299_1, 
        PHYMON_EN_G4398, SRAM_RDATA_SEL_4, Disconnect_C, BACK_EN5715, 
        SUBSID12936_4, IOBA262401, Disconnect_F4934, DEBUGA3249_6, n_5666, 
        TMOUT_PARM4236_4, PHYOPT33553_0, PHYOPTGH3667_6, n_6202, 
        SRAM_RDATA_SEL_30, SRAM_RDATA_SEL_17, DPE13NX, PHYOPTGH3667_1, 
        IOBA82687, SRAM_RDATA_SEL_10, n_10228, n_6724, IOBA222574, 
        SUBSID12936_3, DEBUGB3287_4, DEBUGF_2, SUBSID1_5, Disconnect_D, 
        SRAM_RDATA_SEL_3, PHYOPT33553_7, n_11538, PHYOPT13477_4, 
        TMOUT_PARM4236_3, DEBUGA3249_1, n_2800, SUBSID0_5, SUBVID12860_0, 
        TERMON_B, PHYOPT43591_0, LAT_TM2299_6, SPAREO7, DEBUG02974_1, 
        DEBUG23050_4, REVID_BACK_3, INTLN2337_0, TERMON_A4503, RxData_C, 
        DPE12NX, n_6718, DEBUGD3363_1, DEBUGE3401_5, SUBVID02822_4, n_6190, 
        SUBSID02898_2, PHYOPTEF3629_3, REVID_BACK5677_6, RxData_F4946, 
        SRAM_RDATA_SEL_19, PHYOPT23515_5, n_8202, PHYMON_EN_B, SRAM_SEL5343_1, 
        DEBUGF3439_5, SLAVEMODE4162, DEBUG13012_4, n_10880, n_5668, 
        DEBUG33088_7, Squelch_C4685, a5192, CFGX0, DEBUGC3325_2, INTLN_3, 
        TERMON_E4843, PHYMON_EN_C4374, SRAM_ADDR_IN_6, SRAM_RDATA_SEL_25, 
        Squelch_G5025, DEBUG83126_3, n_11544, PHYOPT13477_6, CACHLN12170, 
        DEBUGD3363_3, n_10216, RxData_A, DEBUG23050_6, INTLN2337_2, 
        REVID_BACK_1, LAT_TM2299_4, DEBUG02974_3, SRAM_LAT_RDATA, SPAREO5, 
        n_10890, PHYOPT43591_2, SUBSID0_7, SUBVID12860_2, PHYMON_EN_B4368, 
        Disconnect_H5104, PHYOPT33553_5, n_2802, DEBUGA3249_3, 
        TMOUT_PARM4236_1, Disconnect_F, BIST_RUN4051, RxDataDly3781_1, 
        SRAM_RDATA_SEL_1, SUBSID12936_1, PHYMON_EN_A4362, RxData_H5116, TSERRS, 
        DEBUGB3287_6, n_6726, SRAM_RDATA_SEL_12, PHYOPTGH3667_3, TTABORTR, 
        n_11546, IOBA302425, Disconnect_B4594, Squelch_B4600, DEBUG9_0, 
        DEBUG83126_1, SRAM_ADDR_IN_4, SRAM_RDATA_SEL_27, RxData_H, INTLN_1, 
        n_5132, IOBA202562, IOSPACE2034, DEBUGC3325_0, SRAM_RUN_2T, 
        DEBUG33088_5, Squelch_B, n_10882, DEBUG13012_6, SRAM_RDATA_SEL_8, 
        DEBUGF3439_7, PHYOPT23515_7, REVID_BACK5677_4, PHYOPTEF3629_1, 
        IOBA142723, SUBVID02822_6, SUBSID02898_0, n_6192, TEST_EYE_EN4274, 
        DEBUGE3401_7, n_10224, PHYOPTEF3629_6, REVID_BACK5677_3, n_6728, 
        PHYOPT23515_0, RxData_B4606, DEBUGE3401_0, SUBSID02898_7, 
        SUBVID02822_1, Disconnect_A4509, n_8042, n_5140, Disconnect_H, 
        DEBUGF3439_0, PHYMON_EN_G, DEBUG13012_1, Squelch_E, DEBUG33088_2, 
        BIST_ERROR, DEBUGC3325_7, n_9562, DEBUG83126_6, n_10218, LAT_TM_6, 
        CACHLN72206, SRAM_RDATA_SEL_20, SRAM_ADDR_IN_3, SRAM_RDATA_SEL_15, 
        n_9570, n_6200, Disconnect_E4849, PHYOPTGH3667_4, n_5664, 
        TMOUT_PARM4236_6, DEBUGA3249_4, PHYOPT33553_2, DEBUGB3287_1, DEBUGF_7, 
        SUBSID12936_6, SUBSID1_0, SRAM_RDATA_SEL_6, Disconnect_A, SPAREO2, 
        DEBUG02974_4, LAT_TM2299_3, REVID_BACK_6, INTLN2337_5, Squelch_H5110, 
        DEBUG23050_1, n_5658, SUBVID12860_5, n_8050, SUBSID0_0, PHYOPT43591_5, 
        TERMON_G, n_11548, DEBUGD3363_4, PHYOPT13477_1, SRAM_RDATA_SEL_29, 
        RxData_F, LockSpd3705_1, DEBUG83126_7, IOBA212568, SUBVID1_2, n_11540, 
        n_2796, n_5134, n_6732, SRAM_ADDR_IN_2, SRAM_RDATA_SEL_21, Squelch_D, 
        TERMON_G5013, DEBUG33088_3, DEBUGC3325_6, n_10884, DEBUGF3439_1, 
        IOBA152729, PHYMON_EN_F, DEBUG13012_0, PHYOPT23515_1, REVID_BACK5677_2, 
        PHYOPTEF3629_7, IOBA272407, DEBUGE3401_1, SUBSID02898_6, n_6194, 
        SUBVID02822_0, DEBUGD3363_5, PHYOPT13477_0, SRAM_RDATA_SEL_28, 
        RxData_G, LockSpd3705_0, SPAREO3, IOBA192556, DEBUG02974_5, IOBA122711, 
        LAT_TM2299_2, SRAM_WR5337, INTLN2337_4, REVID_BACK_7, DEBUG23050_0, 
        SPAREO1_, SUBVID12860_4, SUBSID0_1, PHYOPT43591_4, CACHLN52194, 
        TERMON_F, DEBUGA3249_5, n_2804, TMOUT_PARM4236_7, PHYOPT33553_3, 
        IOBA172544, DEBUGB3287_0, SUBSID12936_7, SRAM_RDATA_SEL_7, 
        PHYMON_EN_E4386, SRAM_RDATA_SEL_14, PHYMON_EN_H4404, n_6720, n_9556, 
        PHYOPTGH3667_5, SRAM_RDATA_SEL_13, PHYOPTGH3667_2, Disconnect_C4679, 
        FastStart3819, PHYOPT33553_4, CLKOFF_EN3164, n_5662, TMOUT_PARM4236_0, 
        DEBUGA3249_2, Disconnect_G, RxDataDly3781_0, PHYMON_EN_H, 
        SRAM_RDATA_SEL_0, SUBSID12936_0, DEBUGB3287_7, DEBUG23050_7, 
        REVID_BACK_0, INTLN2337_3, LAT_TM2299_5, DEBUG02974_2, SPAREO4, 
        TERMON_A, PHYOPT43591_3, SUBSID0_6, IOBA252395, IOBA92693, 
        SUBVID12860_3, PHYOPT13477_7, DEBUGD3363_2, n_2798, RxData_E4861, 
        Squelch_A4515, n_10230, SLAVE_ACT_T, PHYOPT23515_6, DPE14NX, 
        PHYOPTEF3629_0, REVID_BACK5677_5, n_10222, SUBVID02822_7, 
        SUBSID02898_1, DEBUGE3401_6, n_9558, DEBUG0_0, n_8044, INTLN_0, 
        DEBUG13012_7, PHYMON_EN_A, SRAM_RDATA_SEL_9, DEBUGF3439_6, 
        TERMON_B4588, DEBUGC3325_1, DEBUG33088_4, Squelch_C, n_5670, TERMON_H, 
        n_6188, n_9564, DEBUG83126_0, SRAM_RDATA_SEL_26, SRAM_ADDR_IN_5, 
        LAT_TM_0, Squelch_E4855, RxData_A4521, n6145, n6146, n6337, n6338, 
        n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, 
        n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, 
        n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, 
        n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, 
        n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, 
        n6389, n6390, n6391, n6392, n6393, n6395, n6397, n6398, n6399, n6400, 
        n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, 
        n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, 
        n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, 
        n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, 
        n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, 
        n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, 
        n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, 
        n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, 
        n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, 
        n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, 
        n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, 
        n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, 
        n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, 
        n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, 
        n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, 
        n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, 
        n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, 
        n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, 
        n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, 
        n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, 
        n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, 
        n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, 
        n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, 
        n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, 
        n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, 
        n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, 
        n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, 
        n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, 
        n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, 
        n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, 
        n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, 
        n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, 
        n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, 
        n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, 
        n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, 
        n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, 
        n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, 
        n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, 
        n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, 
        n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, 
        n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, 
        n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, 
        n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, 
        n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, 
        n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, 
        n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, 
        n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, 
        n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, 
        n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, 
        n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, 
        n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, 
        n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, 
        n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, 
        n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, 
        n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, 
        n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, 
        n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, 
        n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, 
        n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, 
        n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, 
        n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, 
        n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, 
        n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, 
        n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, 
        n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, 
        n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, 
        n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, 
        n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, 
        n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, 
        n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, 
        n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, 
        n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, 
        n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, 
        n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140;
    assign PCI1WAIT = 1'b0;
    assign ENTXDLY_1 = 1'b0;
    assign DISTXDLY2 = 1'b0;
    assign DISFFCRC0 = 1'b0;
    assign DISFFCRC1 = 1'b0;
    assign DISPFIFO = 1'b0;
    assign DISPFIFO2 = 1'b0;
    assign DISRXZERO = 1'b0;
    assign ENBMUSMRST = 1'b0;
    assign SLQUEUEADDR[1] = 1'b0;
    assign SLQUEUEADDR[0] = 1'b0;
    zan2b REDNT003 ( .A(FBCYC), .B(FB2BKENR), .Y(FB2BKEN) );
    zdffqrb dpe13 ( .CK(PCICLK_FREE), .D(DPE13NX), .R(HRST_), .Q(TMABORTS) );
    zoai21b SPARE755 ( .A(SPAREO1), .B(SRAM_LAT_RDATA), .C(SPAREO9), .Y(
        SPAREO3) );
    zaoi211b SPARE752 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zdffqrb dpe14 ( .CK(PCICLK), .D(DPE14NX), .R(HRST_), .Q(TSERRS) );
    znd2b REDNT002 ( .A(REVID0), .B(1'b0), .Y(DEVS0) );
    zaoi211b SPARE753 ( .A(SPAREO4), .B(n6356), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zoai21b SPARE754 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zdffqrb dpe12 ( .CK(PCICLK_FREE), .D(DPE12NX), .R(HRST_), .Q(TTABORTR) );
    zivb DNTFB2BKENR ( .A(1'b1), .Y(FB2BKENR) );
    zivb DNTSERREN ( .A(1'b1), .Y(SERREN) );
    znr3b SPARE756 ( .A(SPAREO2), .B(CFGX0), .C(SPAREO0_), .Y(SPAREO4) );
    zdffrb SPARE751 ( .CK(PCICLK), .D(SPAREO7), .R(HRST_), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE758 ( .A(SPAREO5), .Y(SPAREO6) );
    znr2b REDNT001 ( .A(REVID0), .B(1'b1), .Y(FBCYC) );
    zdffrb SPARE750 ( .CK(PCICLK), .D(1'b0), .R(HRST_), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb DNTPTER ( .A(1'b1), .Y(RPTYERR) );
    znd3b SPARE759 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb DNTRSTEP ( .A(1'b1), .Y(RSTEP) );
    zivb SPARE757 ( .A(SPAREO4), .Y(SPAREO5) );
    znr3b U1608 ( .A(SRAM_ADDR_IN_2), .B(SRAM_ADDR_IN_0), .C(SRAM_ADDR_IN_6), 
        .Y(n6404) );
    znr2b U1609 ( .A(SRAM_ADDR_IN_3), .B(SRAM_ADDR_IN_4), .Y(n6406) );
    znr2b U1610 ( .A(SRAM_ADDR_IN_5), .B(SRAM_ADDR_IN_1), .Y(n6405) );
    znd2b U1611 ( .A(n6403), .B(n6409), .Y(n6400) );
    znr2b U1612 ( .A(SRAM_ADDR_IN_7), .B(n6386), .Y(n6403) );
    znd2b U1613 ( .A(n6408), .B(n6407), .Y(n6409) );
    znd2b U1614 ( .A(n6386), .B(n6402), .Y(n6408) );
    znd3b U1615 ( .A(n6405), .B(n6406), .C(n6404), .Y(n6407) );
    zor2b U1616 ( .A(PA5I), .B(PA7I), .Y(n6644) );
    zor2b U1617 ( .A(n6398), .B(n6612), .Y(n6742) );
    zoai21b U1618 ( .A(AD2I), .B(AD1I), .C(AD0I), .Y(n6431) );
    znd2b U1619 ( .A(SRAM_RUN_2T), .B(n6616), .Y(n6615) );
    zor2b U1620 ( .A(n6646), .B(n6879), .Y(n6588) );
    zivb U1621 ( .A(n6646), .Y(n6420) );
    znd2b U1622 ( .A(n6411), .B(n6410), .Y(a5192) );
    znd2b U1623 ( .A(n6401), .B(n6386), .Y(n6411) );
    zivb U1624 ( .A(n6409), .Y(n6401) );
    znd2b U1625 ( .A(SRAM_ADDR_IN_8), .B(n6400), .Y(n6410) );
    zivb U1626 ( .A(PA7I), .Y(n6813) );
    zor2b U1627 ( .A(PA7I), .B(n6606), .Y(n6607) );
    zivb U1628 ( .A(PA5I), .Y(n6606) );
    zan3b U1629 ( .A(BACK_EN), .B(n6602), .C(n6419), .Y(n6601) );
    zao22b U1630 ( .A(CP0), .B(n7070), .C(n6361), .D(SUBVID0_0), .Y(n7113) );
    zao22b U1631 ( .A(USBLEGCTLSTS[1]), .B(n6389), .C(PWR_STATE1), .D(n6362), 
        .Y(n7107) );
    zao22b U1632 ( .A(BIST_PATTERN[1]), .B(n7059), .C(CP1), .D(n7070), .Y(
        n7109) );
    zao21b U1633 ( .A(USBLEGCTLSTS[3]), .B(n7125), .C(n6363), .Y(n7087) );
    zoai2x4b U1634 ( .A(n7132), .B(n6986), .C(n7131), .D(n6962), .E(n7134), 
        .F(n6623), .G(n7137), .H(n6872), .Y(n7081) );
    zor2b U1635 ( .A(REVID_BACK_4), .B(n7025), .Y(n7080) );
    zor2b U1636 ( .A(REVID_BACK_7), .B(n7025), .Y(n7076) );
    zao22b U1637 ( .A(SLQUEUEADDR[8]), .B(n7065), .C(n7066), .D(TERMON_A), .Y(
        n7064) );
    zao22b U1638 ( .A(EN_DBG_PORT), .B(n6593), .C(n7072), .D(SRAM_ADDR[8]), 
        .Y(n7071) );
    zao21b U1639 ( .A(REVID0), .B(n7058), .C(n7037), .Y(n7102) );
    zao22b U1640 ( .A(TXDELAY_PARM[1]), .B(n7063), .C(DEBUGE_1), .D(n6593), 
        .Y(n7101) );
    zan2b U1641 ( .A(ENUSB2), .B(PORTWAKECAP3), .Y(n7098) );
    zor2b U1642 ( .A(n6610), .B(n6611), .Y(n6614) );
    zor2b U1643 ( .A(n6611), .B(n6814), .Y(n6815) );
    zor2b U1644 ( .A(n6729), .B(n6878), .Y(n7024) );
    zivb U1645 ( .A(FUNCSEL[2]), .Y(n7021) );
    zivb U1646 ( .A(FUNCSEL[0]), .Y(n7038) );
    zivb U1647 ( .A(FUNCSEL[1]), .Y(n7039) );
    zan2b U1648 ( .A(ENUSB4), .B(PORTWAKECAP7), .Y(n7093) );
    zor2b U1649 ( .A(n6611), .B(n6700), .Y(n7126) );
    zao21b U1650 ( .A(SRAM_RUN), .B(n7072), .C(n7036), .Y(n7090) );
    zor2b U1651 ( .A(n6610), .B(n6611), .Y(n7134) );
    zor2b U1652 ( .A(n6611), .B(n6645), .Y(n7139) );
    zan2b U1653 ( .A(DEBUGF_2), .B(n6593), .Y(n6594) );
    zor2b U1654 ( .A(n6611), .B(n6645), .Y(n7140) );
    zor2b U1655 ( .A(n7036), .B(n7037), .Y(n7035) );
    zor2b U1656 ( .A(n6701), .B(n6878), .Y(n7026) );
    zan2b U1657 ( .A(DEBUGF_3), .B(n6593), .Y(n6592) );
    zor2b U1658 ( .A(n6700), .B(n6701), .Y(n6702) );
    zor2b U1659 ( .A(n6729), .B(n6766), .Y(n6784) );
    zor2b U1660 ( .A(n6645), .B(n6701), .Y(n7138) );
    zor2b U1661 ( .A(n6631), .B(n6700), .Y(n7128) );
    zor2b U1662 ( .A(n6700), .B(n6729), .Y(n7131) );
    zan2b U1663 ( .A(USBLEGCTLSTS[29]), .B(n6425), .Y(n6591) );
    zor2b U1664 ( .A(n6729), .B(n6825), .Y(n6882) );
    zor2b U1665 ( .A(n6631), .B(n6700), .Y(n7129) );
    zor2b U1666 ( .A(n6610), .B(n6631), .Y(n6635) );
    zor2b U1667 ( .A(n6645), .B(n6701), .Y(n6844) );
    zor2b U1668 ( .A(n6700), .B(n6729), .Y(n6934) );
    zor2b U1669 ( .A(n6611), .B(n6878), .Y(n6879) );
    zor2b U1670 ( .A(n6700), .B(n6701), .Y(n7132) );
    zor2b U1671 ( .A(n6611), .B(n6700), .Y(n7127) );
    zivb U1672 ( .A(n6922), .Y(n7074) );
    zor2b U1673 ( .A(n6610), .B(n6611), .Y(n7135) );
    zor2b U1674 ( .A(n6611), .B(n6645), .Y(n6647) );
    zor2b U1675 ( .A(n6631), .B(n6880), .Y(n6881) );
    zao22b U1676 ( .A(SL_ERROFFSET[7]), .B(n7062), .C(USBLEGSUP[31]), .D(n6422
        ), .Y(n7085) );
    zor2b U1677 ( .A(n6701), .B(n6825), .Y(n6883) );
    zor2b U1678 ( .A(n6631), .B(n6824), .Y(n7031) );
    zivb U1679 ( .A(E_PME_EN), .Y(n7032) );
    zor2b U1680 ( .A(n6645), .B(n6701), .Y(n7137) );
    zor2b U1681 ( .A(n6631), .B(n6700), .Y(n6991) );
    zor2b U1682 ( .A(PA2I), .B(PA3I), .Y(n6631) );
    zivb U1683 ( .A(n6631), .Y(CFGX0) );
    zor2b U1684 ( .A(n6700), .B(n6729), .Y(n7130) );
    zor2b U1685 ( .A(n6700), .B(n6701), .Y(n7133) );
    zor2b U1686 ( .A(PA2I), .B(n6699), .Y(n6701) );
    zor2b U1687 ( .A(n6729), .B(n6766), .Y(n7136) );
    zivb U1688 ( .A(PA4I), .Y(n6609) );
    zor2b U1689 ( .A(n6605), .B(n6699), .Y(n6729) );
    zivb U1690 ( .A(PA3I), .Y(n6699) );
    zivb U1691 ( .A(n6729), .Y(n6602) );
    zor2b U1692 ( .A(n6611), .B(n6700), .Y(n6877) );
    zor2b U1693 ( .A(PA3I), .B(n6605), .Y(n6611) );
    zivb U1694 ( .A(PA2I), .Y(n6605) );
    zivb U1695 ( .A(n6611), .Y(n7075) );
    zmux21lb U1696 ( .A(n6385), .B(n6589), .S(n6379), .Y(SRAM_SEL5343_1) );
    zmux21lb U1697 ( .A(n6801), .B(n6590), .S(n6379), .Y(SRAM_SEL5343_0) );
    zivb U1698 ( .A(n6437), .Y(n7055) );
    zmux21lb U1699 ( .A(n7007), .B(n6691), .S(n6358), .Y(DEBUG13012_7) );
    zmux21lb U1700 ( .A(n7008), .B(n6689), .S(n6358), .Y(DEBUG13012_6) );
    zmux21lb U1701 ( .A(n7009), .B(n6687), .S(n6358), .Y(DEBUG13012_5) );
    zmux21lb U1702 ( .A(n7010), .B(n6685), .S(n6358), .Y(DEBUG13012_4) );
    zmux21lb U1703 ( .A(n7011), .B(n6683), .S(n6358), .Y(DEBUG13012_3) );
    zmux21lb U1704 ( .A(TRAP_OPT), .B(n6681), .S(n6358), .Y(DEBUG13012_2) );
    zmux21lb U1705 ( .A(n7012), .B(n6679), .S(n6358), .Y(DEBUG13012_1) );
    zmux21hb U1706 ( .A(DBGIRQ), .B(AD8I), .S(n6358), .Y(DEBUG13012_0) );
    zmux21lb U1707 ( .A(n6992), .B(n6659), .S(n6344), .Y(DEBUG33088_7) );
    zmux21lb U1708 ( .A(n6993), .B(n6587), .S(n6344), .Y(DEBUG33088_6) );
    zmux21lb U1709 ( .A(n6994), .B(n6589), .S(n6344), .Y(DEBUG33088_5) );
    zmux21lb U1710 ( .A(n6995), .B(n6590), .S(n6344), .Y(DEBUG33088_4) );
    zmux21lb U1711 ( .A(n6996), .B(n6654), .S(n6344), .Y(DEBUG33088_3) );
    zmux21lb U1712 ( .A(n6997), .B(n6652), .S(n6344), .Y(DEBUG33088_2) );
    zmux21lb U1713 ( .A(n6998), .B(n6650), .S(n6344), .Y(DEBUG33088_1) );
    zmux21lb U1714 ( .A(n6999), .B(n6648), .S(n6344), .Y(DEBUG33088_0) );
    zmux21lb U1715 ( .A(n6975), .B(n6676), .S(n6352), .Y(DEBUGA3249_7) );
    zmux21lb U1716 ( .A(n6976), .B(n6674), .S(n6352), .Y(DEBUGA3249_6) );
    zmux21lb U1717 ( .A(n6977), .B(n6672), .S(n6352), .Y(DEBUGA3249_5) );
    zmux21lb U1718 ( .A(n6978), .B(n6670), .S(n6352), .Y(DEBUGA3249_4) );
    zmux21lb U1719 ( .A(n6979), .B(n6668), .S(n6352), .Y(DEBUGA3249_3) );
    zmux21lb U1720 ( .A(n6980), .B(n6666), .S(n6352), .Y(DEBUGA3249_2) );
    zmux21lb U1721 ( .A(n6981), .B(n6664), .S(n6352), .Y(DEBUGA3249_1) );
    zmux21lb U1722 ( .A(n6982), .B(n6662), .S(n6352), .Y(DEBUGA3249_0) );
    zmux21lb U1723 ( .A(n6943), .B(n6676), .S(n6338), .Y(DEBUGE3401_7) );
    zmux21lb U1724 ( .A(n6944), .B(n6674), .S(n6338), .Y(DEBUGE3401_6) );
    zmux21lb U1725 ( .A(n6945), .B(n6672), .S(n6338), .Y(DEBUGE3401_5) );
    zmux21lb U1726 ( .A(n6946), .B(n6670), .S(n6338), .Y(DEBUGE3401_4) );
    zmux21lb U1727 ( .A(n6947), .B(n6668), .S(n6338), .Y(DEBUGE3401_3) );
    zmux21lb U1728 ( .A(n6948), .B(n6666), .S(n6338), .Y(DEBUGE3401_2) );
    zmux21lb U1729 ( .A(n6949), .B(n6664), .S(n6338), .Y(DEBUGE3401_1) );
    zmux21lb U1730 ( .A(n6950), .B(n6662), .S(n6338), .Y(DEBUGE3401_0) );
    zmux21lb U1731 ( .A(n6935), .B(n6659), .S(n6350), .Y(DEBUGF3439_7) );
    zmux21lb U1732 ( .A(n6936), .B(n6587), .S(n6350), .Y(DEBUGF3439_6) );
    zmux21lb U1733 ( .A(n6937), .B(n6589), .S(n6350), .Y(DEBUGF3439_5) );
    zmux21lb U1734 ( .A(n6938), .B(n6590), .S(n6350), .Y(DEBUGF3439_4) );
    zmux21lb U1735 ( .A(n6939), .B(n6654), .S(n6350), .Y(DEBUGF3439_3) );
    zmux21lb U1736 ( .A(n6940), .B(n6652), .S(n6350), .Y(DEBUGF3439_2) );
    zmux21lb U1737 ( .A(n6941), .B(n6650), .S(n6350), .Y(DEBUGF3439_1) );
    zmux21lb U1738 ( .A(n6942), .B(n6648), .S(n6350), .Y(DEBUGF3439_0) );
    zmux21lb U1739 ( .A(n6816), .B(n6691), .S(n6349), .Y(REVID_BACK5677_7) );
    zmux21lb U1740 ( .A(n6817), .B(n6689), .S(n6349), .Y(REVID_BACK5677_6) );
    zmux21lb U1741 ( .A(n6818), .B(n6687), .S(n6349), .Y(REVID_BACK5677_5) );
    zmux21lb U1742 ( .A(n6819), .B(n6685), .S(n6349), .Y(REVID_BACK5677_4) );
    zmux21lb U1743 ( .A(n6820), .B(n6683), .S(n6349), .Y(REVID_BACK5677_3) );
    zmux21lb U1744 ( .A(n6821), .B(n6681), .S(n6349), .Y(REVID_BACK5677_2) );
    zmux21lb U1745 ( .A(n6822), .B(n6679), .S(n6349), .Y(REVID_BACK5677_1) );
    zmux21lb U1746 ( .A(n6823), .B(n6634), .S(n6349), .Y(REVID_BACK5677_0) );
    zmux21lb U1747 ( .A(n6791), .B(n6650), .S(n6377), .Y(SUBSID12936_1) );
    zmux21lb U1748 ( .A(n6912), .B(n6666), .S(n6384), .Y(IOBA182550) );
    zmux21hb U1749 ( .A(Squelch_H), .B(SquelchOut_H), .S(PHYMON_EN_H), .Y(
        Squelch_H5110) );
    zmux21lb U1750 ( .A(n6708), .B(n6689), .S(n6341), .Y(n_2798) );
    zmux21lb U1751 ( .A(n6853), .B(n6676), .S(n6343), .Y(PHYOPT33553_7) );
    zmux21lb U1752 ( .A(n6663), .B(n6662), .S(n6355), .Y(n_6202) );
    zmux21lb U1753 ( .A(n6905), .B(n6650), .S(n6383), .Y(IOBA252395) );
    zmux21lb U1754 ( .A(n6897), .B(n6679), .S(n6382), .Y(IOBA92693) );
    zmux41b U1755 ( .A(n6397), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[16]), .D1(
        SRAM_RDATA2[16]), .D2(SRAM_RDATA3[16]), .D3(SRAM_RDATA4[16]), .Y(
        SRAM_RDATA_SEL_16) );
    zmux21lb U1756 ( .A(n7003), .B(n6668), .S(n6340), .Y(DEBUG23050_3) );
    zmux21lb U1757 ( .A(n6834), .B(n6664), .S(n6345), .Y(PHYOPTGH3667_1) );
    zmux21hb U1758 ( .A(TERMON_B), .B(TERM_ON_B), .S(PHYMON_EN_B), .Y(
        TERMON_B4588) );
    zmux21lb U1759 ( .A(n6861), .B(n6691), .S(n6347), .Y(PHYOPT23515_7) );
    zmux41b U1760 ( .A(n6145), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[1]), .D1(
        SRAM_RDATA2[1]), .D2(SRAM_RDATA3[1]), .D3(SRAM_RDATA4[1]), .Y(
        SRAM_RDATA_SEL_1) );
    zmux21lb U1761 ( .A(n6846), .B(n6587), .S(n6359), .Y(PHYOPT43591_6) );
    zmux21lb U1762 ( .A(n6899), .B(n6659), .S(n6383), .Y(IOBA312431) );
    zmux21lb U1763 ( .A(n6843), .B(n6634), .S(n6339), .Y(PHYOPTEF3629_0) );
    zmux21lb U1764 ( .A(n6737), .B(n6683), .S(n6357), .Y(TMOUT_PARM4236_3) );
    zmux21hb U1765 ( .A(Squelch_F), .B(SquelchOut_F), .S(PHYMON_EN_F), .Y(
        Squelch_F4940) );
    zmux41b U1766 ( .A(SRAM_SEL[0]), .B(n6395), .D0(SRAM_RDATA1[23]), .D1(
        SRAM_RDATA2[23]), .D2(SRAM_RDATA3[23]), .D3(SRAM_RDATA4[23]), .Y(
        SRAM_RDATA_SEL_23) );
    zmux21lb U1767 ( .A(n6914), .B(n6662), .S(n6384), .Y(IOBA162538) );
    zmux21lb U1768 ( .A(n6677), .B(n6676), .S(n6355), .Y(n_6188) );
    zmux21lb U1769 ( .A(n6970), .B(n6590), .S(n7053), .Y(DEBUGB3287_4) );
    zmux21lb U1770 ( .A(n6771), .B(n6685), .S(n6375), .Y(SUBVID12860_4) );
    zmux41b U1771 ( .A(n6397), .B(n6395), .D0(SRAM_RDATA1[27]), .D1(
        SRAM_RDATA2[27]), .D2(SRAM_RDATA3[27]), .D3(SRAM_RDATA4[27]), .Y(
        SRAM_RDATA_SEL_27) );
    zmux21lb U1772 ( .A(n6655), .B(n6654), .S(n6351), .Y(n_6726) );
    zmux21lb U1773 ( .A(n6893), .B(n6681), .S(n6346), .Y(LAT_TM2299_2) );
    zmux21lb U1774 ( .A(n6953), .B(n6687), .S(n6354), .Y(DEBUGD3363_5) );
    zmux21lb U1775 ( .A(n6799), .B(n6664), .S(n6378), .Y(SUBSID02898_1) );
    zmux21lb U1776 ( .A(n6745), .B(n6626), .S(n6432), .Y(TEST_EYE_EN4274) );
    zivb U1777 ( .A(AD5I), .Y(n6626) );
    zmux21hb U1778 ( .A(RxData_D), .B(RxDataOut_D), .S(PHYMON_EN_D), .Y(
        RxData_D4776) );
    zmux21lb U1779 ( .A(n6794), .B(n6674), .S(n6378), .Y(SUBSID02898_6) );
    zmux21hb U1780 ( .A(TERMON_H), .B(TERM_ON_H), .S(PHYMON_EN_H), .Y(
        TERMON_H5098) );
    zmux21lb U1781 ( .A(n6772), .B(n6683), .S(n6375), .Y(SUBVID12860_3) );
    zmux21lb U1782 ( .A(n6971), .B(n6654), .S(n7053), .Y(DEBUGB3287_3) );
    zmux21lb U1783 ( .A(n6667), .B(n6666), .S(n6355), .Y(n_6198) );
    zmux41b U1784 ( .A(SRAM_SEL[0]), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[18]), 
        .D1(SRAM_RDATA2[18]), .D2(SRAM_RDATA3[18]), .D3(SRAM_RDATA4[18]), .Y(
        SRAM_RDATA_SEL_18) );
    zmux21lb U1785 ( .A(n6956), .B(n6681), .S(n6354), .Y(DEBUGD3363_2) );
    zmux21lb U1786 ( .A(n6890), .B(n6687), .S(n6346), .Y(LAT_TM2299_5) );
    zmux41b U1787 ( .A(SRAM_SEL[0]), .B(n6395), .D0(SRAM_RDATA1[8]), .D1(
        SRAM_RDATA2[8]), .D2(SRAM_RDATA3[8]), .D3(SRAM_RDATA4[8]), .Y(
        SRAM_RDATA_SEL_8) );
    zmux21lb U1788 ( .A(n6924), .B(n6628), .S(n6432), .Y(FORCE_CRCERR4311) );
    zivb U1789 ( .A(AD6I), .Y(n6628) );
    znd2b U1790 ( .A(HCHALT), .B(n6744), .Y(n6743) );
    zivb U1791 ( .A(n6742), .Y(n6744) );
    zmux21lb U1792 ( .A(n6918), .B(n6685), .S(n6382), .Y(IOBA122711) );
    zmux21lb U1793 ( .A(n6836), .B(n6691), .S(n6339), .Y(PHYOPTEF3629_7) );
    zmux21lb U1794 ( .A(n6736), .B(n6685), .S(n6357), .Y(TMOUT_PARM4236_4) );
    zmux21hb U1795 ( .A(Squelch_B), .B(SquelchOut_B), .S(PHYMON_EN_B), .Y(
        Squelch_B4600) );
    zmux21lb U1796 ( .A(n6868), .B(n6634), .S(n6347), .Y(PHYOPT23515_0) );
    zmux41b U1797 ( .A(n6397), .B(n6395), .D0(SRAM_RDATA1[6]), .D1(SRAM_RDATA2
        [6]), .D2(SRAM_RDATA3[6]), .D3(SRAM_RDATA4[6]), .Y(SRAM_RDATA_SEL_6)
         );
    zmux21lb U1798 ( .A(n6851), .B(n6650), .S(n6359), .Y(PHYOPT43591_1) );
    zmux21hb U1799 ( .A(TERMON_F), .B(TERM_ON_F), .S(PHYMON_EN_F), .Y(
        TERMON_F4928) );
    zmux21lb U1800 ( .A(n6767), .B(n6670), .S(n6340), .Y(DEBUG23050_4) );
    zmux21lb U1801 ( .A(n6829), .B(n6674), .S(n6345), .Y(PHYOPTGH3667_6) );
    znd2b U1802 ( .A(SRAM_ADDR_IN_1), .B(n6637), .Y(n6638) );
    zmux21lb U1803 ( .A(n6860), .B(n6662), .S(n6343), .Y(PHYOPT33553_0) );
    zmux41b U1804 ( .A(n6397), .B(n6395), .D0(SRAM_RDATA1[29]), .D1(
        SRAM_RDATA2[29]), .D2(SRAM_RDATA3[29]), .D3(SRAM_RDATA4[29]), .Y(
        SRAM_RDATA_SEL_29) );
    zmux21lb U1805 ( .A(n6657), .B(n6589), .S(n6351), .Y(n_6722) );
    zmux21lb U1806 ( .A(n6909), .B(n6672), .S(n6384), .Y(IOBA212568) );
    zmux21lb U1807 ( .A(n6786), .B(n6587), .S(n6377), .Y(SUBSID12936_6) );
    zmux21lb U1808 ( .A(n6704), .B(n6679), .S(n6341), .Y(n_2806) );
    zmux41b U1809 ( .A(n6397), .B(n6395), .D0(SRAM_RDATA1[10]), .D1(
        SRAM_RDATA2[10]), .D2(SRAM_RDATA3[10]), .D3(SRAM_RDATA4[10]), .Y(
        SRAM_RDATA_SEL_10) );
    zmux21hb U1810 ( .A(Disconnect_D), .B(DisconnectOut_D), .S(PHYMON_EN_D), 
        .Y(Disconnect_D4764) );
    zmux21lb U1811 ( .A(n6682), .B(n6681), .S(n6337), .Y(n_5668) );
    zmux21lb U1812 ( .A(n6916), .B(n6689), .S(n6382), .Y(IOBA142723) );
    zmux41b U1813 ( .A(SRAM_SEL[0]), .B(n6395), .D0(SRAM_RDATA1[7]), .D1(
        SRAM_RDATA2[7]), .D2(SRAM_RDATA3[7]), .D3(SRAM_RDATA4[7]), .Y(
        SRAM_RDATA_SEL_7) );
    zmux21lb U1814 ( .A(n6867), .B(n6679), .S(n6347), .Y(PHYOPT23515_1) );
    zmux21hb U1815 ( .A(Squelch_D), .B(SquelchOut_D), .S(PHYMON_EN_D), .Y(
        Squelch_D4770) );
    zmux21lb U1816 ( .A(n6852), .B(n6648), .S(n6359), .Y(PHYOPT43591_0) );
    zmux21lb U1817 ( .A(n6837), .B(n6689), .S(n6339), .Y(PHYOPTEF3629_6) );
    zmux21lb U1818 ( .A(n6735), .B(n6687), .S(n6357), .Y(TMOUT_PARM4236_5) );
    zmux21lb U1819 ( .A(n6773), .B(n6681), .S(n6375), .Y(SUBVID12860_2) );
    zmux21lb U1820 ( .A(n6972), .B(n6652), .S(n7053), .Y(DEBUGB3287_2) );
    zmux21lb U1821 ( .A(n6669), .B(n6668), .S(n6355), .Y(n_6196) );
    zmux21hb U1822 ( .A(RxData_B), .B(RxDataOut_B), .S(PHYMON_EN_B), .Y(
        RxData_B4606) );
    zmux41b U1823 ( .A(n6397), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[19]), .D1(
        SRAM_RDATA2[19]), .D2(SRAM_RDATA3[19]), .D3(SRAM_RDATA4[19]), .Y(
        SRAM_RDATA_SEL_19) );
    zmux41b U1824 ( .A(SRAM_SEL[0]), .B(n6395), .D0(SRAM_RDATA1[9]), .D1(
        SRAM_RDATA2[9]), .D2(SRAM_RDATA3[9]), .D3(SRAM_RDATA4[9]), .Y(
        SRAM_RDATA_SEL_9) );
    zmux21lb U1825 ( .A(n6891), .B(n6685), .S(n6346), .Y(LAT_TM2299_4) );
    zmux21lb U1826 ( .A(n6955), .B(n6683), .S(n6354), .Y(DEBUGD3363_3) );
    zmux21lb U1827 ( .A(n6901), .B(n6589), .S(n6383), .Y(IOBA292419) );
    zmux21lb U1828 ( .A(n6793), .B(n6676), .S(n6378), .Y(SUBSID02898_7) );
    zmux41b U1829 ( .A(SRAM_SEL[0]), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[11]), 
        .D1(SRAM_RDATA2[11]), .D2(SRAM_RDATA3[11]), .D3(SRAM_RDATA4[11]), .Y(
        SRAM_RDATA_SEL_11) );
    zmux21lb U1830 ( .A(n6684), .B(n6683), .S(n6337), .Y(n_5666) );
    zmux21hb U1831 ( .A(Disconnect_B), .B(DisconnectOut_B), .S(PHYMON_EN_B), 
        .Y(Disconnect_B4594) );
    zmux21lb U1832 ( .A(n6785), .B(n6659), .S(n6377), .Y(SUBSID12936_7) );
    zmux21lb U1833 ( .A(n6703), .B(n6634), .S(n6341), .Y(n_2808) );
    zmux21lb U1834 ( .A(n6859), .B(n6664), .S(n6343), .Y(PHYOPT33553_1) );
    zmux21lb U1835 ( .A(n6656), .B(n6590), .S(n6351), .Y(n_6724) );
    zmux41b U1836 ( .A(n6397), .B(n6395), .D0(SRAM_RDATA1[28]), .D1(
        SRAM_RDATA2[28]), .D2(SRAM_RDATA3[28]), .D3(SRAM_RDATA4[28]), .Y(
        SRAM_RDATA_SEL_28) );
    zan2b U1837 ( .A(n6379), .B(AD25I), .Y(SRAM_RUN5389) );
    zmux21lb U1838 ( .A(n7002), .B(n6672), .S(n6340), .Y(DEBUG23050_5) );
    zmux21lb U1839 ( .A(n6903), .B(n6654), .S(n6383), .Y(IOBA272407) );
    zmux21lb U1840 ( .A(n6828), .B(n6676), .S(n6345), .Y(PHYOPTGH3667_7) );
    zmux21lb U1841 ( .A(n6907), .B(n6676), .S(n6384), .Y(IOBA232580) );
    zmux21lb U1842 ( .A(n7004), .B(n6666), .S(n6340), .Y(DEBUG23050_2) );
    zmux21lb U1843 ( .A(n6835), .B(n6662), .S(n6345), .Y(PHYOPTGH3667_0) );
    zmux21lb U1844 ( .A(n6854), .B(n6674), .S(n6343), .Y(PHYOPT33553_6) );
    zmux21lb U1845 ( .A(n6665), .B(n6664), .S(n6355), .Y(n_6200) );
    zmux41b U1846 ( .A(n6397), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[17]), .D1(
        SRAM_RDATA2[17]), .D2(SRAM_RDATA3[17]), .D3(SRAM_RDATA4[17]), .Y(
        SRAM_RDATA_SEL_17) );
    zmux21hb U1847 ( .A(TERMON_D), .B(TERM_ON_D), .S(PHYMON_EN_D), .Y(
        TERMON_D4758) );
    zmux21hb U1848 ( .A(RxData_H), .B(RxDataOut_H), .S(PHYMON_EN_H), .Y(
        RxData_H5116) );
    zmux21lb U1849 ( .A(n6792), .B(n6648), .S(n6377), .Y(SUBSID12936_0) );
    zmux21hb U1850 ( .A(Disconnect_F), .B(DisconnectOut_F), .S(PHYMON_EN_F), 
        .Y(Disconnect_F4934) );
    zmux21lb U1851 ( .A(n6603), .B(n6634), .S(n6583), .Y(n_8202) );
    zan2b U1852 ( .A(n6433), .B(n6584), .Y(n6583) );
    zivb U1853 ( .A(n6610), .Y(n6584) );
    zmux21lb U1854 ( .A(n6709), .B(n6691), .S(n6341), .Y(n_2796) );
    zmux21lb U1855 ( .A(n6800), .B(n6662), .S(n6378), .Y(SUBSID02898_0) );
    zmux21lb U1856 ( .A(n6969), .B(n6589), .S(n7053), .Y(DEBUGB3287_5) );
    zmux21lb U1857 ( .A(n6770), .B(n6687), .S(n6375), .Y(SUBVID12860_5) );
    zmux21hb U1858 ( .A(RxData_F), .B(RxDataOut_F), .S(PHYMON_EN_F), .Y(
        RxData_F4946) );
    zmux41b U1859 ( .A(n6397), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[26]), .D1(
        SRAM_RDATA2[26]), .D2(SRAM_RDATA3[26]), .D3(SRAM_RDATA4[26]), .Y(
        SRAM_RDATA_SEL_26) );
    zmux21lb U1860 ( .A(n6653), .B(n6652), .S(n6351), .Y(n_6728) );
    zmux21lb U1861 ( .A(n6892), .B(n6683), .S(n6346), .Y(LAT_TM2299_3) );
    zmux21lb U1862 ( .A(n6954), .B(n6685), .S(n6354), .Y(DEBUGD3363_4) );
    zmux21hb U1863 ( .A(Disconnect_H), .B(DisconnectOut_H), .S(PHYMON_EN_H), 
        .Y(Disconnect_H5104) );
    zmux21lb U1864 ( .A(n6842), .B(n6679), .S(n6339), .Y(PHYOPTEF3629_1) );
    zmux21lb U1865 ( .A(n6738), .B(n6681), .S(n6357), .Y(TMOUT_PARM4236_2) );
    zmux41b U1866 ( .A(SRAM_SEL[0]), .B(n6395), .D0(SRAM_RDATA1[22]), .D1(
        SRAM_RDATA2[22]), .D2(SRAM_RDATA3[22]), .D3(SRAM_RDATA4[22]), .Y(
        SRAM_RDATA_SEL_22) );
    zmux21lb U1867 ( .A(n6675), .B(n6674), .S(n6355), .Y(n_6190) );
    zmux21lb U1868 ( .A(n6862), .B(n6689), .S(n6347), .Y(PHYOPT23515_6) );
    zmux41b U1869 ( .A(n6145), .B(n6146), .D0(SRAM_RDATA1[0]), .D1(SRAM_RDATA2
        [0]), .D2(SRAM_RDATA3[0]), .D3(SRAM_RDATA4[0]), .Y(SRAM_RDATA_SEL_0)
         );
    zmux21lb U1870 ( .A(n6845), .B(n6659), .S(n6359), .Y(PHYOPT43591_7) );
    zmux21lb U1871 ( .A(n6920), .B(n6681), .S(n6382), .Y(IOBA102699) );
    zmux41b U1872 ( .A(n6397), .B(n6395), .D0(SRAM_RDATA1[14]), .D1(
        SRAM_RDATA2[14]), .D2(SRAM_RDATA3[14]), .D3(SRAM_RDATA4[14]), .Y(
        SRAM_RDATA_SEL_14) );
    zmux21lb U1873 ( .A(n6690), .B(n6689), .S(n6337), .Y(n_5660) );
    zmux21hb U1874 ( .A(Squelch_E), .B(SquelchOut_E), .S(PHYMON_EN_E), .Y(
        Squelch_E4855) );
    zmux21lb U1875 ( .A(n6915), .B(n6691), .S(n6382), .Y(IOBA152729) );
    zmux21lb U1876 ( .A(n6790), .B(n6652), .S(n6377), .Y(SUBSID12936_2) );
    zmux21lb U1877 ( .A(n6902), .B(n6590), .S(n6383), .Y(IOBA282413) );
    zmux21lb U1878 ( .A(n6856), .B(n6670), .S(n6343), .Y(PHYOPT33553_4) );
    zmux21lb U1879 ( .A(n6833), .B(n6666), .S(n6345), .Y(PHYOPTGH3667_2) );
    zmux21lb U1880 ( .A(n7006), .B(n6662), .S(n6340), .Y(DEBUG23050_0) );
    zivb U1881 ( .A(AD16I), .Y(n6662) );
    zmux21hb U1882 ( .A(RxData_C), .B(RxDataOut_C), .S(PHYMON_EN_C), .Y(
        RxData_C4691) );
    zmux21lb U1883 ( .A(n6921), .B(n6681), .S(n6380), .Y(INTR_DIS2113) );
    zmux21lb U1884 ( .A(n6847), .B(n6589), .S(n6359), .Y(PHYOPT43591_5) );
    zmux21hb U1885 ( .A(Disconnect_C), .B(DisconnectOut_C), .S(PHYMON_EN_C), 
        .Y(Disconnect_C4679) );
    zmux21lb U1886 ( .A(n6864), .B(n6685), .S(n6347), .Y(PHYOPT23515_4) );
    zmux21lb U1887 ( .A(n6678), .B(n6634), .S(n6337), .Y(n_5672) );
    zmux41b U1888 ( .A(n6145), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[2]), .D1(
        SRAM_RDATA2[2]), .D2(SRAM_RDATA3[2]), .D3(SRAM_RDATA4[2]), .Y(
        SRAM_RDATA_SEL_2) );
    zmux21lb U1889 ( .A(n6671), .B(n6670), .S(n6355), .Y(n_6194) );
    zmux41b U1890 ( .A(SRAM_SEL[0]), .B(n6395), .D0(SRAM_RDATA1[20]), .D1(
        SRAM_RDATA2[20]), .D2(SRAM_RDATA3[20]), .D3(SRAM_RDATA4[20]), .Y(
        SRAM_RDATA_SEL_20) );
    zmux21lb U1891 ( .A(n6840), .B(n6683), .S(n6339), .Y(PHYOPTEF3629_3) );
    zmux21lb U1892 ( .A(n6740), .B(n6634), .S(n6357), .Y(TMOUT_PARM4236_0) );
    zmux21lb U1893 ( .A(n6649), .B(n6648), .S(n6351), .Y(n_6732) );
    zmux21lb U1894 ( .A(n6894), .B(n6679), .S(n6346), .Y(LAT_TM2299_1) );
    zmux21lb U1895 ( .A(n6952), .B(n6689), .S(n6354), .Y(DEBUGD3363_6) );
    zmux21lb U1896 ( .A(n6904), .B(n6652), .S(n6383), .Y(IOBA262401) );
    zmux41b U1897 ( .A(SRAM_SEL[0]), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[24]), 
        .D1(SRAM_RDATA2[24]), .D2(SRAM_RDATA3[24]), .D3(SRAM_RDATA4[24]), .Y(
        SRAM_RDATA_SEL_24) );
    zmux21lb U1898 ( .A(n6967), .B(n6659), .S(n7053), .Y(DEBUGB3287_7) );
    zmux21lb U1899 ( .A(n6768), .B(n6691), .S(n6375), .Y(SUBVID12860_7) );
    zmux21lb U1900 ( .A(n7048), .B(n6618), .S(n6428), .Y(SLAVEMODE4162) );
    zao21b U1901 ( .A(SLAVE_ACT_T), .B(n7044), .C(n6802), .Y(n7048) );
    zivb U1902 ( .A(n6743), .Y(n6432) );
    zmux21lb U1903 ( .A(n6798), .B(n6666), .S(n6378), .Y(SUBSID02898_2) );
    zmux21hb U1904 ( .A(TERMON_A), .B(TERM_ON_A), .S(PHYMON_EN_A), .Y(
        TERMON_A4503) );
    zmux21hb U1905 ( .A(TERMON_E), .B(TERM_ON_E), .S(PHYMON_EN_E), .Y(
        TERMON_E4843) );
    zmux21lb U1906 ( .A(n6795), .B(n6672), .S(n6378), .Y(SUBSID02898_5) );
    zmux21lb U1907 ( .A(n6957), .B(n6679), .S(n6354), .Y(DEBUGD3363_1) );
    zmux21lb U1908 ( .A(n6889), .B(n6689), .S(n6346), .Y(LAT_TM2299_6) );
    zmux21lb U1909 ( .A(n6908), .B(n6674), .S(n6384), .Y(IOBA222574) );
    zmux21lb U1910 ( .A(n6775), .B(n6634), .S(n6375), .Y(SUBVID12860_0) );
    zmux21lb U1911 ( .A(n6974), .B(n6648), .S(n7053), .Y(DEBUGB3287_0) );
    zor2b U1912 ( .A(n6646), .B(n6702), .Y(n7115) );
    zivb U1913 ( .A(n6814), .Y(n6419) );
    zmux21lb U1914 ( .A(n6839), .B(n6685), .S(n6339), .Y(PHYOPTEF3629_4) );
    zmux21lb U1915 ( .A(n6733), .B(n6691), .S(n6357), .Y(TMOUT_PARM4236_7) );
    zmux21lb U1916 ( .A(n6616), .B(n6648), .S(n6379), .Y(SRAM_WR5337) );
    zmux21lb U1917 ( .A(n6850), .B(n6652), .S(n6359), .Y(PHYOPT43591_2) );
    zivb U1918 ( .A(AD26I), .Y(n6652) );
    zmux21hb U1919 ( .A(Disconnect_G), .B(DisconnectOut_G), .S(PHYMON_EN_G), 
        .Y(Disconnect_G5019) );
    zmux41b U1920 ( .A(n6397), .B(n6395), .D0(SRAM_RDATA1[5]), .D1(SRAM_RDATA2
        [5]), .D2(SRAM_RDATA3[5]), .D3(SRAM_RDATA4[5]), .Y(SRAM_RDATA_SEL_5)
         );
    zmux21lb U1921 ( .A(n6865), .B(n6683), .S(n6347), .Y(PHYOPT23515_3) );
    zmux21lb U1922 ( .A(n6830), .B(n6672), .S(n6345), .Y(PHYOPTGH3667_5) );
    zmux21hb U1923 ( .A(RxData_G), .B(RxDataOut_G), .S(PHYMON_EN_G), .Y(
        RxData_G5031) );
    zmux21lb U1924 ( .A(n7000), .B(n6676), .S(n6340), .Y(DEBUG23050_7) );
    zivb U1925 ( .A(AD23I), .Y(n6676) );
    zmux21lb U1926 ( .A(n6857), .B(n6668), .S(n6343), .Y(PHYOPT33553_3) );
    zmux21lb U1927 ( .A(n6919), .B(n6683), .S(n6382), .Y(IOBA112705) );
    zmux21lb U1928 ( .A(n6705), .B(n6681), .S(n6341), .Y(n_2804) );
    zmux41b U1929 ( .A(SRAM_SEL[0]), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[31]), 
        .D1(SRAM_RDATA2[31]), .D2(SRAM_RDATA3[31]), .D3(SRAM_RDATA4[31]), .Y(
        SRAM_RDATA_SEL_31) );
    zmux21lb U1930 ( .A(n6787), .B(n6589), .S(n6377), .Y(SUBSID12936_5) );
    zmux21hb U1931 ( .A(Squelch_A), .B(SquelchOut_A), .S(PHYMON_EN_A), .Y(
        Squelch_A4515) );
    zmux21lb U1932 ( .A(n6660), .B(n6659), .S(n6351), .Y(n_6718) );
    zivb U1933 ( .A(AD31I), .Y(n6659) );
    zmux21lb U1934 ( .A(n6688), .B(n6687), .S(n6337), .Y(n_5662) );
    zivc U1935 ( .A(AD0I), .Y(n6618) );
    zmux41b U1936 ( .A(SRAM_SEL[0]), .B(n6395), .D0(SRAM_RDATA1[13]), .D1(
        SRAM_RDATA2[13]), .D2(SRAM_RDATA3[13]), .D3(SRAM_RDATA4[13]), .Y(
        SRAM_RDATA_SEL_13) );
    zmux21lb U1937 ( .A(n6849), .B(n6654), .S(n6359), .Y(PHYOPT43591_3) );
    zmux41b U1938 ( .A(SRAM_SEL[0]), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[4]), 
        .D1(SRAM_RDATA2[4]), .D2(SRAM_RDATA3[4]), .D3(SRAM_RDATA4[4]), .Y(
        SRAM_RDATA_SEL_4) );
    zmux21lb U1939 ( .A(n6911), .B(n6668), .S(n6384), .Y(IOBA192556) );
    zmux21lb U1940 ( .A(n6866), .B(n6681), .S(n6347), .Y(PHYOPT23515_2) );
    zmux21hb U1941 ( .A(Disconnect_A), .B(DisconnectOut_A), .S(PHYMON_EN_A), 
        .Y(Disconnect_A4509) );
    zmux21lb U1942 ( .A(n6838), .B(n6687), .S(n6339), .Y(PHYOPTEF3629_5) );
    zmux21lb U1943 ( .A(n6734), .B(n6689), .S(n6357), .Y(TMOUT_PARM4236_6) );
    zmux21hb U1944 ( .A(TERMON_C), .B(TERM_ON_C), .S(PHYMON_EN_C), .Y(
        TERMON_C4673) );
    zmux21lb U1945 ( .A(n6888), .B(n6691), .S(n6346), .Y(LAT_TM2299_7) );
    zmux21lb U1946 ( .A(n6958), .B(n6634), .S(n6354), .Y(DEBUGD3363_0) );
    zmux21lb U1947 ( .A(n6774), .B(n6679), .S(n6375), .Y(SUBVID12860_1) );
    zmux21lb U1948 ( .A(n6973), .B(n6650), .S(n7053), .Y(DEBUGB3287_1) );
    zivc U1949 ( .A(n7115), .Y(n7053) );
    zmux21lb U1950 ( .A(n6906), .B(n6648), .S(n6383), .Y(IOBA242389) );
    zivb U1951 ( .A(AD24I), .Y(n6648) );
    zmux21lb U1952 ( .A(n6796), .B(n6670), .S(n6378), .Y(SUBSID02898_4) );
    zmux21lb U1953 ( .A(n6898), .B(n6634), .S(n6382), .Y(IOBA82687) );
    zmux21lb U1954 ( .A(n6900), .B(n6587), .S(n6383), .Y(IOBA302425) );
    zmux21lb U1955 ( .A(n6913), .B(n6664), .S(n6384), .Y(IOBA172544) );
    zmux21lb U1956 ( .A(n6686), .B(n6685), .S(n6337), .Y(n_5664) );
    zmux21hb U1957 ( .A(Squelch_G), .B(SquelchOut_G), .S(PHYMON_EN_G), .Y(
        Squelch_G5025) );
    zmux41b U1958 ( .A(SRAM_SEL[0]), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[12]), 
        .D1(SRAM_RDATA2[12]), .D2(SRAM_RDATA3[12]), .D3(SRAM_RDATA4[12]), .Y(
        SRAM_RDATA_SEL_12) );
    zmux21lb U1959 ( .A(n6706), .B(n6683), .S(n6341), .Y(n_2802) );
    zivb U1960 ( .A(AD11I), .Y(n6683) );
    zmux41b U1961 ( .A(n6397), .B(n6395), .D0(SRAM_RDATA1[30]), .D1(
        SRAM_RDATA2[30]), .D2(SRAM_RDATA3[30]), .D3(SRAM_RDATA4[30]), .Y(
        SRAM_RDATA_SEL_30) );
    zmux21lb U1962 ( .A(n6788), .B(n6590), .S(n6377), .Y(SUBSID12936_4) );
    zmux21lb U1963 ( .A(n6658), .B(n6587), .S(n6351), .Y(n_6720) );
    zmux21hb U1964 ( .A(RxData_A), .B(RxDataOut_A), .S(PHYMON_EN_A), .Y(
        RxData_A4521) );
    zmux21lb U1965 ( .A(n6858), .B(n6666), .S(n6343), .Y(PHYOPT33553_2) );
    zivb U1966 ( .A(AD18I), .Y(n6666) );
    zmux21lb U1967 ( .A(n6831), .B(n6670), .S(n6345), .Y(PHYOPTGH3667_4) );
    zmux21lb U1968 ( .A(n7001), .B(n6674), .S(n6340), .Y(DEBUG23050_6) );
    zivb U1969 ( .A(AD22I), .Y(n6674) );
    zmux21lb U1970 ( .A(n6832), .B(n6668), .S(n6345), .Y(PHYOPTGH3667_3) );
    zmux21lb U1971 ( .A(n7005), .B(n6664), .S(n6340), .Y(DEBUG23050_1) );
    zivb U1972 ( .A(AD17I), .Y(n6664) );
    zmux21lb U1973 ( .A(n6855), .B(n6672), .S(n6343), .Y(PHYOPT33553_5) );
    zmux21hb U1974 ( .A(RxData_E), .B(RxDataOut_E), .S(PHYMON_EN_E), .Y(
        RxData_E4861) );
    zmux21lb U1975 ( .A(n7020), .B(n6687), .S(n6341), .Y(CLKOFF_EN3164) );
    znr2b U1976 ( .A(n6632), .B(n7133), .Y(n6341) );
    zmux21lb U1977 ( .A(n6707), .B(n6685), .S(n6341), .Y(n_2800) );
    zivb U1978 ( .A(AD12I), .Y(n6685) );
    zmux21lb U1979 ( .A(n6789), .B(n6654), .S(n6377), .Y(SUBSID12936_3) );
    zivb U1980 ( .A(AD27I), .Y(n6654) );
    zmux21hb U1981 ( .A(Squelch_C), .B(SquelchOut_C), .S(PHYMON_EN_C), .Y(
        Squelch_C4685) );
    zmux41b U1982 ( .A(SRAM_SEL[0]), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[15]), 
        .D1(SRAM_RDATA2[15]), .D2(SRAM_RDATA3[15]), .D3(SRAM_RDATA4[15]), .Y(
        SRAM_RDATA_SEL_15) );
    zmux21lb U1983 ( .A(n6917), .B(n6687), .S(n6382), .Y(IOBA132717) );
    zmux21lb U1984 ( .A(n6692), .B(n6691), .S(n6337), .Y(n_5658) );
    zmux21lb U1985 ( .A(n6910), .B(n6670), .S(n6384), .Y(IOBA202562) );
    zivb U1986 ( .A(AD20I), .Y(n6670) );
    zmux21lb U1987 ( .A(n6797), .B(n6668), .S(n6378), .Y(SUBSID02898_3) );
    zivb U1988 ( .A(AD19I), .Y(n6668) );
    zmux21lb U1989 ( .A(n6651), .B(n6650), .S(n6351), .Y(n_6730) );
    zivb U1990 ( .A(AD25I), .Y(n6650) );
    zmux21lb U1991 ( .A(n6951), .B(n6691), .S(n6354), .Y(DEBUGD3363_7) );
    zivb U1992 ( .A(AD15I), .Y(n6691) );
    zmux21lb U1993 ( .A(n6895), .B(n6634), .S(n6346), .Y(LAT_TM2299_0) );
    zivb U1994 ( .A(AD8I), .Y(n6634) );
    zmux41b U1995 ( .A(n6397), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[25]), .D1(
        SRAM_RDATA2[25]), .D2(SRAM_RDATA3[25]), .D3(SRAM_RDATA4[25]), .Y(
        SRAM_RDATA_SEL_25) );
    zmux21lb U1996 ( .A(n6769), .B(n6689), .S(n6375), .Y(SUBVID12860_6) );
    zivb U1997 ( .A(AD14I), .Y(n6689) );
    zmux21lb U1998 ( .A(n6968), .B(n6587), .S(n7053), .Y(DEBUGB3287_6) );
    zmux21lb U1999 ( .A(n6430), .B(n6619), .S(n6356), .Y(SWDBG4088) );
    zivb U2000 ( .A(AD1I), .Y(n6619) );
    zmux21hb U2001 ( .A(TERMON_G), .B(TERM_ON_G), .S(PHYMON_EN_G), .Y(
        TERMON_G5013) );
    zmux21lb U2002 ( .A(n6673), .B(n6672), .S(n6355), .Y(n_6192) );
    zivb U2003 ( .A(AD21I), .Y(n6672) );
    zmux41b U2004 ( .A(n6397), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[21]), .D1(
        SRAM_RDATA2[21]), .D2(SRAM_RDATA3[21]), .D3(SRAM_RDATA4[21]), .Y(
        SRAM_RDATA_SEL_21) );
    zmux21hb U2005 ( .A(Disconnect_E), .B(DisconnectOut_E), .S(PHYMON_EN_E), 
        .Y(Disconnect_E4849) );
    zmux21lb U2006 ( .A(n6841), .B(n6681), .S(n6339), .Y(PHYOPTEF3629_2) );
    zivb U2007 ( .A(AD10I), .Y(n6681) );
    zmux21lb U2008 ( .A(n6739), .B(n6679), .S(n6357), .Y(TMOUT_PARM4236_1) );
    zmux21lb U2009 ( .A(n6848), .B(n6590), .S(n6359), .Y(PHYOPT43591_4) );
    zmux21lb U2010 ( .A(n6680), .B(n6679), .S(n6337), .Y(n_5670) );
    zivb U2011 ( .A(AD9I), .Y(n6679) );
    zmux21lb U2012 ( .A(n6863), .B(n6687), .S(n6347), .Y(PHYOPT23515_5) );
    zivb U2013 ( .A(AD13I), .Y(n6687) );
    zmux41b U2014 ( .A(n6397), .B(SRAM_SEL[1]), .D0(SRAM_RDATA1[3]), .D1(
        SRAM_RDATA2[3]), .D2(SRAM_RDATA3[3]), .D3(SRAM_RDATA4[3]), .Y(
        SRAM_RDATA_SEL_3) );
    zivf U2015 ( .A(n6617), .Y(n6436) );
    zivb U2016 ( .A(n6615), .Y(SRAM_LAT_RDATA) );
    zor2b U2017 ( .A(n6413), .B(TABORTR), .Y(DPE12NX) );
    zivb U2018 ( .A(AD28I), .Y(n6590) );
    zor2b U2019 ( .A(n6412), .B(SERRS), .Y(DPE14NX) );
    zivb U2020 ( .A(AD30I), .Y(n6587) );
    zor2b U2021 ( .A(n6423), .B(MABORTS), .Y(DPE13NX) );
    zivb U2022 ( .A(AD29I), .Y(n6589) );
    zivb U2023 ( .A(n6636), .Y(SRAM_ADDR[0]) );
    znd2b U2024 ( .A(SRAM_ADDR_IN_0), .B(n6637), .Y(n6636) );
    zivb U2025 ( .A(n6639), .Y(SRAM_ADDR[2]) );
    znd2b U2026 ( .A(SRAM_ADDR_IN_2), .B(n6637), .Y(n6639) );
    zivb U2027 ( .A(n6640), .Y(SRAM_ADDR[3]) );
    znd2b U2028 ( .A(SRAM_ADDR_IN_3), .B(n6637), .Y(n6640) );
    zivb U2029 ( .A(n6641), .Y(SRAM_ADDR[4]) );
    znd2b U2030 ( .A(SRAM_ADDR_IN_4), .B(n6637), .Y(n6641) );
    zivb U2031 ( .A(n6642), .Y(SRAM_ADDR[5]) );
    znd2b U2032 ( .A(SRAM_ADDR_IN_5), .B(n6637), .Y(n6642) );
    zivb U2033 ( .A(n6643), .Y(SRAM_ADDR[6]) );
    znd2b U2034 ( .A(SRAM_ADDR_IN_6), .B(n6637), .Y(n6643) );
    zivb U2035 ( .A(a5192), .Y(n6637) );
    zivb U2036 ( .A(n6604), .Y(SRAM_ADDR[7]) );
    zmux21lb U2037 ( .A(SRAM_ADDR_IN_7), .B(n6395), .S(a5192), .Y(n6604) );
    zivb U2038 ( .A(n6603), .Y(SRAM_ADDR[8]) );
    zmux21lb U2039 ( .A(SRAM_ADDR_IN_8), .B(n6385), .S(a5192), .Y(n6603) );
    zor2b U2040 ( .A(n6381), .B(n6380), .Y(PCI_RPCMD) );
    zan2b U2041 ( .A(n6586), .B(n6399), .Y(n6424) );
    zan2b U2042 ( .A(n6414), .B(n6427), .Y(PCI_R6DG) );
    zivb U2043 ( .A(n6765), .Y(n6427) );
    zor2b U2044 ( .A(n6632), .B(n6729), .Y(n6765) );
    zan2b U2045 ( .A(n6414), .B(n6415), .Y(PCI_R6CG) );
    zivb U2046 ( .A(n6730), .Y(n6415) );
    zan2b U2047 ( .A(n6362), .B(n6399), .Y(R84G) );
    zan2b U2048 ( .A(n6414), .B(n6433), .Y(R61G) );
    zivb U2049 ( .A(n6825), .Y(n6414) );
    zivb U2050 ( .A(PA6I), .Y(n6608) );
    zivb U2051 ( .A(n6633), .Y(n6433) );
    zor2b U2052 ( .A(n6631), .B(n6632), .Y(n6633) );
    zan2b U2053 ( .A(INTLN_0), .B(n6421), .Y(UIRQSEL0) );
    zan2b U2054 ( .A(INTLN_1), .B(n6421), .Y(UIRQSEL1) );
    zan2b U2055 ( .A(INTLN_2), .B(n6421), .Y(UIRQSEL2) );
    zan2b U2056 ( .A(INTLN_3), .B(n6421), .Y(UIRQSEL3) );
    zao22b U2057 ( .A(SQSET[0]), .B(n6593), .C(BIST_PATTERN[0]), .D(n7059), 
        .Y(n6439) );
    zoai2x4b U2058 ( .A(n6728), .B(n7023), .C(n6756), .D(n7126), .E(n6741), 
        .F(n7044), .G(n6635), .H(n6636), .Y(n6440) );
    zivb U2059 ( .A(SLAVE_ACT), .Y(n7044) );
    zivb U2060 ( .A(n6638), .Y(SRAM_ADDR[1]) );
    zivb U2061 ( .A(n6635), .Y(n7072) );
    zao22b U2062 ( .A(MMSPACE), .B(n7083), .C(SQSET[1]), .D(n6593), .Y(n6443)
         );
    zoai2x4b U2063 ( .A(n6727), .B(n7023), .C(FCFG), .D(n7128), .E(n6754), .F(
        n7126), .G(n6741), .H(n6430), .Y(n6444) );
    zoai2x4b U2064 ( .A(n6726), .B(n7023), .C(n6752), .D(n7127), .E(n6741), 
        .F(n6429), .G(n6635), .H(n6639), .Y(n6446) );
    zao22b U2065 ( .A(BMASTREN), .B(n7083), .C(EN_UTM_RESET), .D(n7063), .Y(
        n6447) );
    zoai2x4b U2066 ( .A(n6781), .B(n6784), .C(n6991), .D(n7018), .E(n6647), 
        .F(n6693), .G(n7024), .H(n7040), .Y(n6451) );
    zoai2x4b U2067 ( .A(n6702), .B(n6987), .C(n7130), .D(n6963), .E(n6614), 
        .F(n6621), .G(n7138), .H(n6873), .Y(n6452) );
    zoai2x4b U2068 ( .A(n6725), .B(n7023), .C(n6750), .D(n7126), .E(n6741), 
        .F(n7034), .G(n6635), .H(n6640), .Y(n6453) );
    zoai2x4b U2069 ( .A(n6780), .B(n7136), .C(n7129), .D(n7017), .E(n6647), 
        .F(n6694), .G(n7024), .H(n7033), .Y(n6455) );
    zoai2x4b U2070 ( .A(n7130), .B(n6961), .C(n7135), .D(n6625), .E(n7137), 
        .F(n6871), .G(n6778), .H(n6784), .Y(n6460) );
    zoai2x4b U2071 ( .A(n6724), .B(n7023), .C(n6748), .D(n7127), .E(n6635), 
        .F(n6642), .G(n6702), .H(n6985), .Y(n6461) );
    zoai2x4b U2072 ( .A(n7131), .B(n6960), .C(n6614), .D(n6627), .E(n7138), 
        .F(n6870), .G(n6777), .H(n7136), .Y(n6464) );
    zoai2x4b U2073 ( .A(n6722), .B(n7023), .C(n6747), .D(n6877), .E(n6635), 
        .F(n6643), .G(n7132), .H(n6984), .Y(n6465) );
    zoai2x4b U2074 ( .A(n6934), .B(n6959), .C(n7134), .D(n6629), .E(n6844), 
        .F(n6869), .G(n6776), .H(n6784), .Y(n6468) );
    zoai2x4b U2075 ( .A(n6723), .B(n7023), .C(n6746), .D(n7126), .E(n6604), 
        .F(n6635), .G(n7133), .H(n6983), .Y(n6469) );
    zoai2x4b U2076 ( .A(n6991), .B(n7012), .C(n6934), .D(n6957), .E(n6894), 
        .F(n7024), .G(n7138), .H(n6867), .Y(n6477) );
    zoai2x4b U2077 ( .A(n6739), .B(n6741), .C(n7133), .D(n6704), .E(n6815), 
        .F(n6822), .G(n6614), .H(n6717), .Y(n6479) );
    zoai2x4b U2078 ( .A(n6879), .B(n6921), .C(n6893), .D(n7024), .E(n7131), 
        .F(n6956), .G(TRAP_OPT), .H(n6991), .Y(n6482) );
    zoai2x4b U2079 ( .A(n6738), .B(n6741), .C(n6702), .D(n6705), .E(n6815), 
        .F(n6821), .G(n7135), .H(n6718), .Y(n6485) );
    zoai2x4b U2080 ( .A(n6772), .B(n6784), .C(n6737), .D(n6741), .E(n7133), 
        .F(n6706), .G(n6815), .H(n6820), .Y(n6488) );
    zoai2x4b U2081 ( .A(n6958), .B(n7031), .C(n7128), .D(n7011), .E(n7130), 
        .F(n6955), .G(n6892), .H(n7024), .Y(n6490) );
    zoai2x4b U2082 ( .A(n6991), .B(n7010), .C(n7130), .D(n6954), .E(n6891), 
        .F(n7024), .G(n6844), .H(n6864), .Y(n6492) );
    zoai2x4b U2083 ( .A(n6736), .B(n6741), .C(n7132), .D(n6707), .E(n6815), 
        .F(n6819), .G(n6614), .H(n6719), .Y(n6494) );
    zoai2x4b U2084 ( .A(n7128), .B(n7009), .C(n7131), .D(n6953), .E(n6890), 
        .F(n7024), .G(n6702), .H(n7020), .Y(n6496) );
    zivb U2085 ( .A(n7026), .Y(n7037) );
    zoai2x4b U2086 ( .A(n6877), .B(n6929), .C(n6735), .D(n6741), .E(n6815), 
        .F(n6818), .G(n7134), .H(n6720), .Y(n6498) );
    zivb U2087 ( .A(n7024), .Y(n7068) );
    zoai2x4b U2088 ( .A(n6763), .B(n6877), .C(n6734), .D(n6741), .E(n6702), 
        .F(n6708), .G(n6815), .H(n6817), .Y(n6502) );
    zao22b U2089 ( .A(USBLEGCTLSTS[15]), .B(n7125), .C(PME_STS), .D(n6362), 
        .Y(n6504) );
    zoai2x4b U2090 ( .A(n6808), .B(n7126), .C(n6733), .D(n6741), .E(n7132), 
        .F(n6709), .G(n6815), .H(n6816), .Y(n6505) );
    zoai2x4b U2091 ( .A(n6958), .B(n7031), .C(n7129), .D(n7007), .E(n6934), 
        .F(n6951), .G(n6888), .H(n7024), .Y(n6507) );
    zoai2x4b U2092 ( .A(n6647), .B(n6663), .C(n6881), .D(n6914), .E(n6753), 
        .F(n7127), .G(n7135), .H(n6712), .Y(n6508) );
    zoai2x4b U2093 ( .A(n7138), .B(n6860), .C(n7133), .D(n6982), .E(n7130), 
        .F(n6950), .G(n7129), .H(n7006), .Y(n6509) );
    zoai2x4b U2094 ( .A(n7129), .B(n7005), .C(n6647), .D(n6665), .E(n6881), 
        .F(n6913), .G(n7127), .H(n6928), .Y(n6512) );
    zoai2x4b U2095 ( .A(n7139), .B(n6667), .C(n6881), .D(n6912), .E(n6762), 
        .F(n6877), .G(n6614), .H(n6713), .Y(n6519) );
    zoai2x4b U2096 ( .A(n6844), .B(n6858), .C(n6702), .D(n6980), .E(n7131), 
        .F(n6948), .G(n6991), .H(n7004), .Y(n6520) );
    zao22b U2097 ( .A(DISPFUNDRN), .B(n7060), .C(SLQUEUEADDR[19]), .D(n7065), 
        .Y(n6522) );
    zoai2x4b U2098 ( .A(E_PME_EN), .B(n7031), .C(n7137), .D(n6857), .E(n7133), 
        .F(n6979), .G(n7131), .H(n6947), .Y(n6523) );
    zoai2x4b U2099 ( .A(n6934), .B(n6946), .C(n7139), .D(n6671), .E(n6881), 
        .F(n6910), .G(n7134), .H(n6714), .Y(n6530) );
    zoai2x4b U2100 ( .A(n6767), .B(n6991), .C(n7138), .D(n6856), .E(n6751), 
        .F(n7126), .G(n7132), .H(n6978), .Y(n6531) );
    zoai2x4b U2101 ( .A(n6991), .B(n7002), .C(n7140), .D(n6673), .E(n6881), 
        .F(n6909), .G(n7135), .H(n6715), .Y(n6535) );
    zoai2x4b U2102 ( .A(n6844), .B(n6855), .C(n7126), .D(n6927), .E(n6702), 
        .F(n6977), .G(n7130), .H(n6945), .Y(n6536) );
    zivb U2103 ( .A(n6815), .Y(n7058) );
    zoai2x4b U2104 ( .A(n7128), .B(n7001), .C(n6647), .D(n6675), .E(n6881), 
        .F(n6908), .G(n6614), .H(n6716), .Y(n6540) );
    zoai2x4b U2105 ( .A(n7137), .B(n6854), .C(n6761), .D(n6877), .E(n7132), 
        .F(n6976), .G(n6934), .H(n6944), .Y(n6541) );
    zao222b U2106 ( .A(BIST_PATTERN[23]), .B(n7059), .C(IOBA23), .D(n6586), 
        .E(CTRL_G[3]), .F(n7069), .Y(n6542) );
    zao22b U2107 ( .A(SELEOF), .B(n7060), .C(SLQUEUEADDR[23]), .D(n7065), .Y(
        n6543) );
    zoai2x4b U2108 ( .A(n7138), .B(n6853), .C(n6807), .D(n7126), .E(n7133), 
        .F(n6975), .G(n7130), .H(n6943), .Y(n6544) );
    zoai2x4b U2109 ( .A(n6635), .B(n6616), .C(n7128), .D(n6999), .E(n6934), 
        .F(n6942), .G(n7137), .H(n6852), .Y(n6548) );
    zoai2x4b U2110 ( .A(n7136), .B(n6791), .C(n7132), .D(n6973), .E(n6881), 
        .F(n6905), .G(n6877), .H(n6926), .Y(n6551) );
    zivb U2111 ( .A(n6879), .Y(n7083) );
    zoai2x4b U2112 ( .A(n6881), .B(n6904), .C(n6760), .D(n7127), .E(n7139), 
        .F(n6653), .G(n7134), .H(n6710), .Y(n6558) );
    zoai2x4b U2113 ( .A(n6881), .B(n6903), .C(n6806), .D(n6877), .E(n7140), 
        .F(n6655), .G(n7135), .H(n6711), .Y(n6562) );
    zao22b U2114 ( .A(CTRL_A[0]), .B(n7070), .C(n7066), .D(TERMON_F), .Y(n6564
        ) );
    zoai2x4b U2115 ( .A(n6879), .B(n6933), .C(n6635), .D(n6801), .E(n7131), 
        .F(n6938), .G(n7128), .H(n6995), .Y(n6565) );
    zivb U2116 ( .A(TTABORTR), .Y(n6933) );
    zivb U2117 ( .A(n7132), .Y(n7063) );
    zao22b U2118 ( .A(CTRL_A[1]), .B(n7070), .C(Disconnect_F), .D(n7066), .Y(
        n6570) );
    zivb U2119 ( .A(n7127), .Y(n7066) );
    zoai2x4b U2120 ( .A(n6879), .B(n6932), .C(n6385), .D(n6635), .E(n7130), 
        .F(n6937), .G(n7129), .H(n6994), .Y(n6571) );
    zivb U2121 ( .A(TMABORTS), .Y(n6932) );
    zao22b U2122 ( .A(IOBA29), .B(n6586), .C(SLQUEUEADDR[29]), .D(n7065), .Y(
        n6573) );
    zoai2x4b U2123 ( .A(n6879), .B(n6931), .C(n6991), .D(n6993), .E(n6934), 
        .F(n6936), .G(n6844), .H(n6846), .Y(n6576) );
    zivb U2124 ( .A(TSERRS), .Y(n6931) );
    zivb U2125 ( .A(n7031), .Y(n7036) );
    zivb U2126 ( .A(n7130), .Y(n6593) );
    zivb U2127 ( .A(n6991), .Y(n7060) );
    zivb U2128 ( .A(n7137), .Y(n7070) );
    zivb U2129 ( .A(n6881), .Y(n6586) );
    zivb U2130 ( .A(n6647), .Y(n7065) );
    zivb U2131 ( .A(n7135), .Y(n7059) );
    zdffrb INTLN_reg_7 ( .CK(PCICLK), .D(INTLN2337_7), .R(HRST_), .QN(n6723)
         );
    zdffrb INTLN_reg_6 ( .CK(PCICLK), .D(INTLN2337_6), .R(HRST_), .QN(n6722)
         );
    zdffrb INTLN_reg_5 ( .CK(PCICLK), .D(INTLN2337_5), .R(HRST_), .QN(n6724)
         );
    zdffrb INTLN_reg_4 ( .CK(PCICLK), .D(INTLN2337_4), .R(HRST_), .Q(INTLN_4), 
        .QN(n6721) );
    zdffqrb INTLN_reg_3 ( .CK(PCICLK), .D(INTLN2337_3), .R(HRST_), .Q(INTLN_3)
         );
    zivb U2132 ( .A(INTLN_3), .Y(n6725) );
    zdffqrb INTLN_reg_2 ( .CK(PCICLK), .D(INTLN2337_2), .R(HRST_), .Q(INTLN_2)
         );
    zivb U2133 ( .A(INTLN_2), .Y(n6726) );
    zdffqrb INTLN_reg_1 ( .CK(PCICLK), .D(INTLN2337_1), .R(HRST_), .Q(INTLN_1)
         );
    zivb U2134 ( .A(INTLN_1), .Y(n6727) );
    zdffqrb INTLN_reg_0 ( .CK(PCICLK), .D(INTLN2337_0), .R(HRST_), .Q(INTLN_0)
         );
    zivb U2135 ( .A(INTLN_0), .Y(n6728) );
    zdffrb DEBUG0_reg_7 ( .CK(PCICLK), .D(DEBUG02974_7), .R(HRST_), .Q(CAHCFG_
        ), .QN(n7013) );
    zdffrb DEBUG0_reg_6 ( .CK(PCICLK), .D(DEBUG02974_6), .R(HRST_), .Q(BABOPT), 
        .QN(n7014) );
    zdffrb DEBUG0_reg_5 ( .CK(PCICLK), .D(DEBUG02974_5), .R(HRST_), .Q(PAROPT), 
        .QN(n7015) );
    zdffrb DEBUG0_reg_4 ( .CK(PCICLK), .D(DEBUG02974_4), .R(HRST_), .Q(REDUCE), 
        .QN(n7016) );
    zdffrb DEBUG0_reg_3 ( .CK(PCICLK), .D(DEBUG02974_3), .R(HRST_), .Q(
        HCISPEC_), .QN(n7017) );
    zdffqrb DEBUG0_reg_2 ( .CK(PCICLK), .D(DEBUG02974_2), .R(HRST_), .Q(PM_EN)
         );
    zivb U2136 ( .A(PM_EN), .Y(n7018) );
    zdffrb DEBUG0_reg_1 ( .CK(PCICLK), .D(DEBUG02974_1), .R(HRST_), .QN(FCFG)
         );
    zdffrb DEBUG0_reg_0 ( .CK(PCICLK), .D(DEBUG02974_0), .R(HRST_), .Q(
        DEBUG0_0), .QN(n7019) );
    zdffrb DEBUG1_reg_7 ( .CK(PCICLK), .D(DEBUG13012_7), .R(HRST_), .Q(
        DISSTUFF), .QN(n7007) );
    zdffrb DEBUG1_reg_6 ( .CK(PCICLK), .D(DEBUG13012_6), .R(HRST_), .Q(DISPRST
        ), .QN(n7008) );
    zdffrb DEBUG1_reg_5 ( .CK(PCICLK), .D(DEBUG13012_5), .R(HRST_), .Q(DISEOP), 
        .QN(n7009) );
    zdffrb DEBUG1_reg_4 ( .CK(PCICLK), .D(DEBUG13012_4), .R(HRST_), .Q(ENOCPY), 
        .QN(n7010) );
    zdffrb DEBUG1_reg_3 ( .CK(PCICLK), .D(DEBUG13012_3), .R(HRST_), .Q(TESTCNT
        ), .QN(n7011) );
    zdffrb DEBUG1_reg_2 ( .CK(PCICLK), .D(DEBUG13012_2), .R(HRST_), .QN(
        TRAP_OPT) );
    zdffrb DEBUG1_reg_1 ( .CK(PCICLK), .D(DEBUG13012_1), .R(HRST_), .Q(VIAPSS), 
        .QN(n7012) );
    zdffqrb DEBUG1_reg_0 ( .CK(PCICLK), .D(DEBUG13012_0), .R(HRST_), .Q(DBGIRQ
        ) );
    zdffrb DEBUG3_reg_7 ( .CK(PCICLK), .D(DEBUG33088_7), .R(HRST_), .Q(
        DIS_TERM_ON_H), .QN(n6992) );
    zdffrb DEBUG3_reg_6 ( .CK(PCICLK), .D(DEBUG33088_6), .R(HRST_), .Q(
        DIS_TERM_ON_G), .QN(n6993) );
    zdffrb DEBUG3_reg_5 ( .CK(PCICLK), .D(DEBUG33088_5), .R(HRST_), .Q(
        DIS_TERM_ON_F), .QN(n6994) );
    zdffrb DEBUG3_reg_4 ( .CK(PCICLK), .D(DEBUG33088_4), .R(HRST_), .Q(
        DIS_TERM_ON_E), .QN(n6995) );
    zdffrb DEBUG3_reg_3 ( .CK(PCICLK), .D(DEBUG33088_3), .R(HRST_), .Q(
        DIS_TERM_ON_D), .QN(n6996) );
    zdffrb DEBUG3_reg_2 ( .CK(PCICLK), .D(DEBUG33088_2), .R(HRST_), .Q(
        DIS_TERM_ON_C), .QN(n6997) );
    zdffrb DEBUG3_reg_1 ( .CK(PCICLK), .D(DEBUG33088_1), .R(HRST_), .Q(
        DIS_TERM_ON_B), .QN(n6998) );
    zdffrb DEBUG3_reg_0 ( .CK(PCICLK), .D(DEBUG33088_0), .R(HRST_), .Q(
        DIS_TERM_ON_A), .QN(n6999) );
    zdffrb DEBUGA_reg_7 ( .CK(PCICLK), .D(DEBUGA3249_7), .R(HRST_), .Q(
        TXDELAY_PARM[7]), .QN(n6975) );
    zdffrb DEBUGA_reg_6 ( .CK(PCICLK), .D(DEBUGA3249_6), .R(HRST_), .Q(
        TXDELAY_PARM[6]), .QN(n6976) );
    zdffrb DEBUGA_reg_5 ( .CK(PCICLK), .D(DEBUGA3249_5), .R(HRST_), .Q(
        TXDELAY_PARM[5]), .QN(n6977) );
    zdffrb DEBUGA_reg_4 ( .CK(PCICLK), .D(DEBUGA3249_4), .R(HRST_), .Q(
        TXDELAY_PARM[4]), .QN(n6978) );
    zdffrb DEBUGA_reg_3 ( .CK(PCICLK), .D(DEBUGA3249_3), .R(HRST_), .Q(
        TXDELAY_PARM[3]), .QN(n6979) );
    zdffrb DEBUGA_reg_2 ( .CK(PCICLK), .D(DEBUGA3249_2), .R(HRST_), .Q(
        TXDELAY_PARM[2]), .QN(n6980) );
    zdffrb DEBUGA_reg_1 ( .CK(PCICLK), .D(DEBUGA3249_1), .R(HRST_), .Q(
        TXDELAY_PARM[1]), .QN(n6981) );
    zdffrb DEBUGA_reg_0 ( .CK(PCICLK), .D(DEBUGA3249_0), .R(HRST_), .Q(
        TXDELAY_PARM[0]), .QN(n6982) );
    zdffrb DEBUGE_reg_7 ( .CK(PCICLK), .D(DEBUGE3401_7), .R(HRST_), .QN(n6943)
         );
    zdffrb DEBUGE_reg_6 ( .CK(PCICLK), .D(DEBUGE3401_6), .R(HRST_), .QN(n6944)
         );
    zdffrb DEBUGE_reg_5 ( .CK(PCICLK), .D(DEBUGE3401_5), .R(HRST_), .QN(n6945)
         );
    zdffrb DEBUGE_reg_4 ( .CK(PCICLK), .D(DEBUGE3401_4), .R(HRST_), .QN(n6946)
         );
    zdffrb DEBUGE_reg_3 ( .CK(PCICLK), .D(DEBUGE3401_3), .R(HRST_), .QN(n6947)
         );
    zdffrb DEBUGE_reg_2 ( .CK(PCICLK), .D(DEBUGE3401_2), .R(HRST_), .QN(n6948)
         );
    zdffrb DEBUGE_reg_1 ( .CK(PCICLK), .D(DEBUGE3401_1), .R(HRST_), .Q(
        DEBUGE_1), .QN(n6949) );
    zdffrb DEBUGE_reg_0 ( .CK(PCICLK), .D(DEBUGE3401_0), .R(HRST_), .QN(n6950)
         );
    zdffrb DEBUGF_reg_7 ( .CK(PCICLK), .D(DEBUGF3439_7), .R(HRST_), .Q(
        DEBUGF_7), .QN(n6935) );
    zdffrb DEBUGF_reg_6 ( .CK(PCICLK), .D(DEBUGF3439_6), .R(HRST_), .QN(n6936)
         );
    zdffrb DEBUGF_reg_5 ( .CK(PCICLK), .D(DEBUGF3439_5), .R(HRST_), .QN(n6937)
         );
    zdffrb DEBUGF_reg_4 ( .CK(PCICLK), .D(DEBUGF3439_4), .R(HRST_), .QN(n6938)
         );
    zdffqrb DEBUGF_reg_3 ( .CK(PCICLK), .D(DEBUGF3439_3), .R(HRST_), .Q(
        DEBUGF_3) );
    zivb U2137 ( .A(DEBUGF_3), .Y(n6939) );
    zdffqrb DEBUGF_reg_2 ( .CK(PCICLK), .D(DEBUGF3439_2), .R(HRST_), .Q(
        DEBUGF_2) );
    zivb U2138 ( .A(DEBUGF_2), .Y(n6940) );
    zdffrb DEBUGF_reg_1 ( .CK(PCICLK), .D(DEBUGF3439_1), .R(HRST_), .QN(n6941)
         );
    zdffrb DEBUGF_reg_0 ( .CK(PCICLK), .D(DEBUGF3439_0), .R(HRST_), .QN(n6942)
         );
    zdffsb LockSpd_reg_1 ( .CK(PCICLK), .D(LockSpd3705_1), .S(HRST_), .Q(
        LockSpd[1]), .QN(n6886) );
    zdffsb LockSpd_reg_0 ( .CK(PCICLK), .D(LockSpd3705_0), .S(HRST_), .Q(
        LockSpd[0]), .QN(n6887) );
    zdffrb TrkSpd_reg_1 ( .CK(PCICLK), .D(TrkSpd3743_1), .R(HRST_), .Q(TrkSpd
        [1]), .QN(n6731) );
    zdffrb TrkSpd_reg_0 ( .CK(PCICLK), .D(TrkSpd3743_0), .R(HRST_), .Q(TrkSpd
        [0]), .QN(n6732) );
    zdffrb REVID_BACK_reg_7 ( .CK(PCICLK), .D(REVID_BACK5677_7), .R(HRST_), 
        .Q(REVID_BACK_7), .QN(n6816) );
    zdffrb REVID_BACK_reg_6 ( .CK(PCICLK), .D(REVID_BACK5677_6), .R(HRST_), 
        .Q(REVID_BACK_6), .QN(n6817) );
    zdffrb REVID_BACK_reg_5 ( .CK(PCICLK), .D(REVID_BACK5677_5), .R(HRST_), 
        .Q(REVID_BACK_5), .QN(n6818) );
    zdffrb REVID_BACK_reg_4 ( .CK(PCICLK), .D(REVID_BACK5677_4), .R(HRST_), 
        .Q(REVID_BACK_4), .QN(n6819) );
    zdffrb REVID_BACK_reg_3 ( .CK(PCICLK), .D(REVID_BACK5677_3), .R(HRST_), 
        .Q(REVID_BACK_3), .QN(n6820) );
    zdffrb REVID_BACK_reg_2 ( .CK(PCICLK), .D(REVID_BACK5677_2), .R(HRST_), 
        .Q(REVID_BACK_2), .QN(n6821) );
    zdffrb REVID_BACK_reg_1 ( .CK(PCICLK), .D(REVID_BACK5677_1), .R(HRST_), 
        .Q(REVID_BACK_1), .QN(n6822) );
    zdffrb REVID_BACK_reg_0 ( .CK(PCICLK), .D(REVID_BACK5677_0), .R(HRST_), 
        .Q(REVID_BACK_0), .QN(n6823) );
    zdffrb SUBVID0_reg_4 ( .CK(PCICLK), .D(SUBVID02822_4), .R(HRST_), .QN(
        n6779) );
    zdffrb DEBUGC_reg_4 ( .CK(PCICLK), .D(DEBUGC3325_4), .R(HRST_), .QN(n6962)
         );
    zdffrb SUBSID1_reg_1 ( .CK(PCICLK), .D(SUBSID12936_1), .R(HRST_), .QN(
        n6791) );
    zdffrb IOBA18_reg ( .CK(PCICLK), .D(IOBA182550), .R(HRST_), .Q(IOBA18), 
        .QN(n6912) );
    zdffqrb SRAM_RUN_2T_reg ( .CK(PCICLK), .D(SRAM_RUN_T), .R(HRST_), .Q(
        SRAM_RUN_2T) );
    zdffrb Squelch_H_reg ( .CK(PCICLK), .D(Squelch_H5110), .R(HRST_), .Q(
        Squelch_H), .QN(n6757) );
    zdffsb DEBUG9_reg_6 ( .CK(PCICLK), .D(n_2798), .S(HRST_), .Q(TXTMOUT_EN), 
        .QN(n6708) );
    zdffsb PHYOPT3_reg_7 ( .CK(PCICLK), .D(PHYOPT33553_7), .S(HRST_), .Q(
        CTRL_C[3]), .QN(n6853) );
    zdffrb SLQUEUE_ADDR_reg3_16 ( .CK(PCICLK), .D(n_6202), .R(HRST_), .Q(
        SLQUEUEADDR[16]), .QN(n6663) );
    zdffrb IOBA25_reg ( .CK(PCICLK), .D(IOBA252395), .R(HRST_), .Q(IOBA25), 
        .QN(n6905) );
    zdffrb CACHLN6_reg ( .CK(PCICLK), .D(CACHLN62200), .R(HRST_), .Q(CACHLN6), 
        .QN(n7028) );
    zdffrb IOBA9_reg ( .CK(PCICLK), .D(IOBA92693), .R(HRST_), .Q(IOBA9), .QN(
        n6897) );
    zdffqrb BIST_PATTERN_reg3_16 ( .CK(PCICLK), .D(n_10890), .R(HRST_), .Q(
        BIST_PATTERN[16]) );
    zivb U2139 ( .A(BIST_PATTERN[16]), .Y(n6712) );
    zdffrb PHYMON_EN_F_reg ( .CK(PCICLK), .D(PHYMON_EN_F4392), .R(HRST_), .Q(
        PHYMON_EN_F), .QN(n6748) );
    zdffrb DEBUG2_reg_3 ( .CK(PCICLK), .D(DEBUG23050_3), .R(HRST_), .Q(
        DISPFUNDRN), .QN(n7003) );
    zdffrb PHYOPTGH_reg_1 ( .CK(PCICLK), .D(PHYOPTGH3667_1), .R(HRST_), .Q(
        CTRL_H[1]), .QN(n6834) );
    zdffrb TERMON_B_reg ( .CK(PCICLK), .D(TERMON_B4588), .R(HRST_), .Q(
        TERMON_B), .QN(n6755) );
    zdffqrb SRAM_ADDR_IN_reg_6 ( .CK(PCICLK), .D(n_8042), .R(HRST_), .Q(
        SRAM_ADDR_IN_6) );
    zdffrb PHYOPT1_reg_3 ( .CK(PCICLK), .D(PHYOPT13477_3), .R(HRST_), .Q(
        loopback), .QN(n6873) );
    zdffrb PHYOPT2_reg_7 ( .CK(PCICLK), .D(PHYOPT23515_7), .R(HRST_), .Q(
        PdPHY_Dis), .QN(n6861) );
    zdffqrb BIST_PATTERN_reg_1 ( .CK(PCICLK), .D(n_9568), .R(HRST_), .Q(
        BIST_PATTERN[1]) );
    zdffsb RxDataDly_reg_2 ( .CK(PCICLK), .D(RxDataDly3781_2), .S(HRST_), .Q(
        RxDataDly[2]), .QN(n6810) );
    zdffrb PHYOPT4_reg_6 ( .CK(PCICLK), .D(PHYOPT43591_6), .R(HRST_), .Q(
        CTRL_A[2]), .QN(n6846) );
    zdffrb IOBA31_reg ( .CK(PCICLK), .D(IOBA312431), .R(HRST_), .Q(IOBA31), 
        .QN(n6899) );
    zdffrb PHYOPTEF_reg_0 ( .CK(PCICLK), .D(PHYOPTEF3629_0), .R(HRST_), .Q(
        CTRL_F[0]), .QN(n6843) );
    zdffrb TMOUT_PARM_reg_3 ( .CK(PCICLK), .D(TMOUT_PARM4236_3), .R(CMDRST_), 
        .Q(TMOUT_PARM[3]), .QN(n6737) );
    zdffrb Squelch_F_reg ( .CK(PCICLK), .D(Squelch_F4940), .R(HRST_), .Q(
        Squelch_F), .QN(n6759) );
    zdffqrb BIST_PATTERN_reg3_23 ( .CK(PCICLK), .D(n_10876), .R(HRST_), .Q(
        BIST_PATTERN[23]) );
    zdffrb IOSPACE_reg ( .CK(PCICLK), .D(IOSPACE2034), .R(HRST_), .Q(IOSPACE), 
        .QN(n6896) );
    zdffrb IOBA16_reg ( .CK(PCICLK), .D(IOBA162538), .R(HRST_), .Q(IOBA16), 
        .QN(n6914) );
    zdffrb SLQUEUE_ADDR_reg3_23 ( .CK(PCICLK), .D(n_6188), .R(HRST_), .Q(
        SLQUEUEADDR[23]), .QN(n6677) );
    zdffrb PHYMON_EN_H_reg ( .CK(PCICLK), .D(PHYMON_EN_H4404), .R(HRST_), .Q(
        PHYMON_EN_H), .QN(n6746) );
    zdffrb DEBUGB_reg_4 ( .CK(PCICLK), .D(DEBUGB3287_4), .R(HRST_), .Q(
        DIS_SOF_RUN), .QN(n6970) );
    zdffsb SUBVID1_reg_4 ( .CK(PCICLK), .D(SUBVID12860_4), .S(HRST_), .QN(
        n6771) );
    zdffqrb BIST_PATTERN_reg4_27 ( .CK(PCICLK), .D(n_11544), .R(HRST_), .Q(
        BIST_PATTERN[27]) );
    zivb U2140 ( .A(BIST_PATTERN[27]), .Y(n6711) );
    zdffrb SLQUEUE_ADDR_reg4_27 ( .CK(PCICLK), .D(n_6726), .R(HRST_), .Q(
        SLQUEUEADDR[27]), .QN(n6655) );
    zdffsb LAT_TM_reg_2 ( .CK(PCICLK), .D(LAT_TM2299_2), .S(HRST_), .QN(n6893)
         );
    zdffrb DEBUGD_reg_5 ( .CK(PCICLK), .D(DEBUGD3363_5), .R(HRST_), .QN(n6953)
         );
    zdffrb SUBSID0_reg_1 ( .CK(PCICLK), .D(SUBSID02898_1), .R(HRST_), .Q(
        SUBSID0_1), .QN(n6799) );
    zdffrb TEST_EYE_EN_reg ( .CK(PCICLK_FREE), .D(TEST_EYE_EN4274), .R(CMDRST_
        ), .Q(TEST_EYE_EN), .QN(n6745) );
    zdffrb DEBUG8_reg_6 ( .CK(PCICLK), .D(DEBUG83126_6), .R(HRST_), .Q(
        ENISOHANDCHK), .QN(n6984) );
    zdffrb RxData_D_reg ( .CK(PCICLK), .D(RxData_D4776), .R(HRST_), .Q(
        RxData_D), .QN(n6807) );
    zdffrb SUBSID0_reg_6 ( .CK(PCICLK), .D(SUBSID02898_6), .R(HRST_), .Q(
        SUBSID0_6), .QN(n6794) );
    zdffsb DEBUG8_reg_1 ( .CK(PCICLK), .D(DEBUG83126_1), .S(HRST_), .Q(
        EN_CHKTOGCRC), .QN(n6989) );
    zdffqrb TERMON_H_reg ( .CK(PCICLK), .D(TERMON_H5098), .R(HRST_), .Q(
        TERMON_H) );
    zdffrb SUBVID1_reg_3 ( .CK(PCICLK), .D(SUBVID12860_3), .R(HRST_), .QN(
        n6772) );
    zdffsb DEBUGB_reg_3 ( .CK(PCICLK), .D(DEBUGB3287_3), .S(HRST_), .Q(
        TURN_PARM[3]), .QN(n6971) );
    zdffrb SLQUEUE_ADDR_reg3_18 ( .CK(PCICLK), .D(n_6198), .R(HRST_), .Q(
        SLQUEUEADDR[18]), .QN(n6667) );
    zdffqrb BIST_PATTERN_reg3_18 ( .CK(PCICLK), .D(n_10886), .R(HRST_), .Q(
        BIST_PATTERN[18]) );
    zivb U2141 ( .A(BIST_PATTERN[18]), .Y(n6713) );
    zdffrb DEBUGD_reg_2 ( .CK(PCICLK), .D(DEBUGD3363_2), .R(HRST_), .QN(n6956)
         );
    zdffrb LAT_TM_reg_5 ( .CK(PCICLK), .D(LAT_TM2299_5), .R(HRST_), .QN(n6890)
         );
    zdffqrb BIST_PATTERN_reg2_8 ( .CK(PCICLK), .D(n_10230), .R(HRST_), .Q(
        BIST_PATTERN[8]) );
    zdffqrb BIST_RUN_reg ( .CK(PCICLK_FREE), .D(BIST_RUN4051), .R(CMDRST_), 
        .Q(BIST_RUN) );
    zivb U2142 ( .A(BIST_RUN), .Y(n6429) );
    zdffrb FORCE_CRCERR_reg ( .CK(PCICLK_FREE), .D(FORCE_CRCERR4311), .R(
        CMDRST_), .Q(FORCE_CRCERR), .QN(n6924) );
    zdffrb IOBA12_reg ( .CK(PCICLK), .D(IOBA122711), .R(HRST_), .Q(IOBA12), 
        .QN(n6918) );
    zdffsb PHYOPTEF_reg_7 ( .CK(PCICLK), .D(PHYOPTEF3629_7), .S(HRST_), .Q(
        CTRL_E[3]), .QN(n6836) );
    zdffrb TMOUT_PARM_reg_4 ( .CK(PCICLK), .D(TMOUT_PARM4236_4), .R(CMDRST_), 
        .Q(TMOUT_PARM[4]), .QN(n6736) );
    zdffrb Squelch_B_reg ( .CK(PCICLK), .D(Squelch_B4600), .R(HRST_), .Q(
        Squelch_B), .QN(n6763) );
    zdffsb PHYOPT2_reg_0 ( .CK(PCICLK), .D(PHYOPT23515_0), .S(HRST_), .Q(
        BypassDiv4), .QN(n6868) );
    zdffqrb BIST_PATTERN_reg_6 ( .CK(PCICLK), .D(n_9558), .R(HRST_), .Q(
        BIST_PATTERN[6]) );
    zivb U2143 ( .A(BIST_PATTERN[6]), .Y(n6627) );
    zdffrb PHYOPT4_reg_1 ( .CK(PCICLK), .D(PHYOPT43591_1), .R(HRST_), .Q(
        CTRL_B[1]), .QN(n6851) );
    zdffqrb TERMON_F_reg ( .CK(PCICLK), .D(TERMON_F4928), .R(HRST_), .Q(
        TERMON_F) );
    zdffrb DEBUG2_reg_4 ( .CK(PCICLK), .D(DEBUG23050_4), .R(HRST_), .Q(SUBIDWE
        ), .QN(n6767) );
    zdffrb PHYOPT1_reg_4 ( .CK(PCICLK), .D(PHYOPT13477_4), .R(HRST_), .Q(
        tstmod), .QN(n6872) );
    zdffrb PHYOPTGH_reg_6 ( .CK(PCICLK), .D(PHYOPTGH3667_6), .R(HRST_), .Q(
        CTRL_G[2]), .QN(n6829) );
    zdffqrb SRAM_ADDR_IN_reg_1 ( .CK(PCICLK), .D(n_8052), .R(HRST_), .Q(
        SRAM_ADDR_IN_1) );
    zdffrb PHYMON_EN_B_reg ( .CK(PCICLK), .D(PHYMON_EN_B4368), .R(HRST_), .Q(
        PHYMON_EN_B), .QN(n6754) );
    zdffrb PHYOPT3_reg_0 ( .CK(PCICLK), .D(PHYOPT33553_0), .R(HRST_), .Q(
        CTRL_D[0]), .QN(n6860) );
    zdffrb CACHLN2_reg ( .CK(PCICLK), .D(CACHLN22176), .R(HRST_), .Q(CACHLN2), 
        .QN(n7040) );
    zdffqrb BIST_PATTERN_reg4_29 ( .CK(PCICLK), .D(n_11540), .R(HRST_), .Q(
        BIST_PATTERN[29]) );
    zdffrb SLQUEUE_ADDR_reg4_29 ( .CK(PCICLK), .D(n_6722), .R(HRST_), .Q(
        SLQUEUEADDR[29]), .QN(n6657) );
    zdffrb IOBA21_reg ( .CK(PCICLK), .D(IOBA212568), .R(HRST_), .Q(IOBA21), 
        .QN(n6909) );
    zdffrb SUBSID1_reg_6 ( .CK(PCICLK), .D(SUBSID12936_6), .R(HRST_), .QN(
        n6786) );
    zdffrb DEBUG9_reg_1 ( .CK(PCICLK), .D(n_2806), .R(HRST_), .QN(n6704) );
    zdffrb SUBVID0_reg_3 ( .CK(PCICLK), .D(SUBVID02822_3), .R(HRST_), .QN(
        n6780) );
    zdffrb DEBUGC_reg_3 ( .CK(PCICLK), .D(DEBUGC3325_3), .R(HRST_), .Q(
        sync_fast), .QN(n6963) );
    zdffrb BIST_ERROR_reg ( .CK(PCICLK_FREE), .D(BIST_ERROR4199), .R(CMDRST_), 
        .Q(BIST_ERROR), .QN(n7034) );
    zdffqrb BIST_PATTERN_reg2_10 ( .CK(PCICLK), .D(n_10226), .R(HRST_), .Q(
        BIST_PATTERN[10]) );
    zivb U2144 ( .A(BIST_PATTERN[10]), .Y(n6718) );
    zdffrb Disconnect_D_reg ( .CK(PCICLK), .D(Disconnect_D4764), .R(HRST_), 
        .Q(Disconnect_D), .QN(n6927) );
    zdffrb SLQUEUE_ADDR_reg2_10 ( .CK(PCICLK), .D(n_5668), .R(HRST_), .Q(
        SLQUEUEADDR[10]), .QN(n6682) );
    zdffrb SLQUEUE_ADDR_reg_6 ( .CK(PCICLK), .D(n_5134), .R(HRST_), .Q(
        SLQUEUEADDR[6]), .QN(n6697) );
    zdffrb IOBA14_reg ( .CK(PCICLK), .D(IOBA142723), .R(HRST_), .Q(IOBA14), 
        .QN(n6916) );
    zdffqrb BIST_PATTERN_reg_7 ( .CK(PCICLK), .D(n_9556), .R(HRST_), .Q(
        BIST_PATTERN[7]) );
    zivb U2145 ( .A(BIST_PATTERN[7]), .Y(n6629) );
    zdffsb PHYOPT2_reg_1 ( .CK(PCICLK), .D(PHYOPT23515_1), .S(HRST_), .Q(TMODE
        ), .QN(n6867) );
    zdffrb Squelch_D_reg ( .CK(PCICLK), .D(Squelch_D4770), .R(HRST_), .Q(
        Squelch_D), .QN(n6761) );
    zdffrb PHYOPT4_reg_0 ( .CK(PCICLK), .D(PHYOPT43591_0), .R(HRST_), .Q(
        CTRL_B[0]), .QN(n6852) );
    zdffrb PHYOPTEF_reg_6 ( .CK(PCICLK), .D(PHYOPTEF3629_6), .R(HRST_), .Q(
        CTRL_E[2]), .QN(n6837) );
    zdffsb TMOUT_PARM_reg_5 ( .CK(PCICLK), .D(TMOUT_PARM4236_5), .S(CMDRST_), 
        .Q(TMOUT_PARM[5]), .QN(n6735) );
    zdffrb SUBVID1_reg_2 ( .CK(PCICLK), .D(SUBVID12860_2), .R(HRST_), .Q(
        SUBVID1_2), .QN(n6773) );
    zdffrb DEBUGB_reg_2 ( .CK(PCICLK), .D(DEBUGB3287_2), .R(HRST_), .Q(
        TURN_PARM[2]), .QN(n6972) );
    zdffrb SLQUEUE_ADDR_reg3_19 ( .CK(PCICLK), .D(n_6196), .R(HRST_), .Q(
        SLQUEUEADDR[19]), .QN(n6669) );
    zdffrb RxData_B_reg ( .CK(PCICLK), .D(RxData_B4606), .R(HRST_), .Q(
        RxData_B), .QN(n6808) );
    zdffqrb BIST_PATTERN_reg3_19 ( .CK(PCICLK), .D(n_10884), .R(HRST_), .Q(
        BIST_PATTERN[19]) );
    zdffqrb BIST_PATTERN_reg2_9 ( .CK(PCICLK), .D(n_10228), .R(HRST_), .Q(
        BIST_PATTERN[9]) );
    zivb U2146 ( .A(BIST_PATTERN[9]), .Y(n6717) );
    zdffsb LAT_TM_reg_4 ( .CK(PCICLK), .D(LAT_TM2299_4), .S(HRST_), .QN(n6891)
         );
    zdffrb DEBUGD_reg_3 ( .CK(PCICLK), .D(DEBUGD3363_3), .R(HRST_), .QN(n6955)
         );
    zdffrb IOBA29_reg ( .CK(PCICLK), .D(IOBA292419), .R(HRST_), .Q(IOBA29), 
        .QN(n6901) );
    zdffrb SUBSID0_reg_7 ( .CK(PCICLK), .D(SUBSID02898_7), .R(HRST_), .Q(
        SUBSID0_7), .QN(n6793) );
    zdffrb DEBUG8_reg_0 ( .CK(PCICLK), .D(DEBUG83126_0), .R(HRST_), .Q(
        HsEnFB_Dis), .QN(n6990) );
    zdffsb SUBVID0_reg_2 ( .CK(PCICLK), .D(SUBVID02822_2), .S(HRST_), .QN(
        n6781) );
    zdffrb DEBUGC_reg_2 ( .CK(PCICLK), .D(DEBUGC3325_2), .R(HRST_), .Q(
        sync_jend), .QN(n6964) );
    zdffqrb BIST_PATTERN_reg2_11 ( .CK(PCICLK), .D(n_10224), .R(HRST_), .Q(
        BIST_PATTERN[11]) );
    zdffrb SLQUEUE_ADDR_reg2_11 ( .CK(PCICLK), .D(n_5666), .R(HRST_), .Q(
        SLQUEUEADDR[11]), .QN(n6684) );
    zdffrb SLQUEUE_ADDR_reg_7 ( .CK(PCICLK), .D(n_5132), .R(HRST_), .Q(
        SLQUEUEADDR[7]), .QN(n6698) );
    zdffrb Disconnect_B_reg ( .CK(PCICLK), .D(Disconnect_B4594), .R(HRST_), 
        .Q(Disconnect_B), .QN(n6929) );
    zdffrb SUBSID1_reg_7 ( .CK(PCICLK), .D(SUBSID12936_7), .R(HRST_), .QN(
        n6785) );
    zdffqrb SRAM_RUN_T_reg ( .CK(PCICLK), .D(SRAM_RUN), .R(HRST_), .Q(
        SRAM_RUN_T) );
    zdffrb DEBUG9_reg_0 ( .CK(PCICLK), .D(n_2808), .R(HRST_), .Q(DEBUG9_0), 
        .QN(n6703) );
    zdffrb PHYOPT3_reg_1 ( .CK(PCICLK), .D(PHYOPT33553_1), .R(HRST_), .Q(
        CTRL_D[1]), .QN(n6859) );
    zdffrb SLQUEUE_ADDR_reg4_28 ( .CK(PCICLK), .D(n_6724), .R(HRST_), .Q(
        SLQUEUEADDR[28]), .QN(n6656) );
    zdffqrb BIST_PATTERN_reg4_28 ( .CK(PCICLK), .D(n_11542), .R(HRST_), .Q(
        BIST_PATTERN[28]) );
    zdffqrb SRAM_RUN_reg ( .CK(PCICLK), .D(SRAM_RUN5389), .R(HRST_), .Q(
        SRAM_RUN) );
    zdffrb PHYMON_EN_D_reg ( .CK(PCICLK), .D(PHYMON_EN_D4380), .R(HRST_), .Q(
        PHYMON_EN_D), .QN(n6750) );
    zdffrb DEBUG2_reg_5 ( .CK(PCICLK), .D(DEBUG23050_5), .R(HRST_), .Q(
        ENTXDLY_2), .QN(n7002) );
    zdffrb CACHLN4_reg ( .CK(PCICLK), .D(CACHLN42188), .R(HRST_), .Q(CACHLN4), 
        .QN(n7030) );
    zdffrb PHYOPT1_reg_5 ( .CK(PCICLK), .D(PHYOPT13477_5), .R(HRST_), .Q(
        rx_block_dis), .QN(n6871) );
    zdffrb IOBA27_reg ( .CK(PCICLK), .D(IOBA272407), .R(HRST_), .Q(IOBA27), 
        .QN(n6903) );
    zdffsb PHYOPTGH_reg_7 ( .CK(PCICLK), .D(PHYOPTGH3667_7), .S(HRST_), .Q(
        CTRL_G[3]), .QN(n6828) );
    zdffqrb SRAM_ADDR_IN_reg_0 ( .CK(PCICLK), .D(n_8054), .R(HRST_), .Q(
        SRAM_ADDR_IN_0) );
    zdffrb IOBA23_reg ( .CK(PCICLK), .D(IOBA232580), .R(HRST_), .Q(IOBA23), 
        .QN(n6907) );
    zdffrb DEBUG2_reg_2 ( .CK(PCICLK), .D(DEBUG23050_2), .R(HRST_), .Q(
        DISTXDLY), .QN(n7004) );
    zdffrb CACHLN0_reg ( .CK(PCICLK), .D(CACHLN02164), .R(HRST_), .Q(CACHLN0), 
        .QN(n7043) );
    zdffsb PHYOPT1_reg_2 ( .CK(PCICLK), .D(PHYOPT13477_2), .S(HRST_), .Q(
        SOF_DISCONN_CHK), .QN(n6874) );
    zdffrb PHYOPTGH_reg_0 ( .CK(PCICLK), .D(PHYOPTGH3667_0), .R(HRST_), .Q(
        CTRL_H[0]), .QN(n6835) );
    zdffrb SRAM_ADDR_IN_reg_7 ( .CK(PCICLK), .D(n_8040), .R(HRST_), .Q(
        SRAM_ADDR_IN_7), .QN(n6402) );
    zdffrb PHYOPT3_reg_6 ( .CK(PCICLK), .D(PHYOPT33553_6), .R(HRST_), .Q(
        CTRL_C[2]), .QN(n6854) );
    zdffrb SLQUEUE_ADDR_reg3_17 ( .CK(PCICLK), .D(n_6200), .R(HRST_), .Q(
        SLQUEUEADDR[17]), .QN(n6665) );
    zdffqrb BIST_PATTERN_reg3_17 ( .CK(PCICLK), .D(n_10888), .R(HRST_), .Q(
        BIST_PATTERN[17]) );
    zdffrb TERMON_D_reg ( .CK(PCICLK), .D(TERMON_D4758), .R(HRST_), .Q(
        TERMON_D), .QN(n6751) );
    zdffrb RxData_H_reg ( .CK(PCICLK), .D(RxData_H5116), .R(HRST_), .Q(
        RxData_H), .QN(n6803) );
    zdffsb SUBSID1_reg_0 ( .CK(PCICLK), .D(SUBSID12936_0), .S(HRST_), .Q(
        SUBSID1_0), .QN(n6792) );
    zdffqrb Disconnect_F_reg ( .CK(PCICLK), .D(Disconnect_F4934), .R(HRST_), 
        .Q(Disconnect_F) );
    zdffqrb SRAM_ADDR_IN_reg2_8 ( .CK(PCICLK), .D(n_8202), .R(HRST_), .Q(
        SRAM_ADDR_IN_8) );
    zdffrb DEBUG9_reg_7 ( .CK(PCICLK), .D(n_2796), .R(HRST_), .Q(TXDELAY_EN), 
        .QN(n6709) );
    zdffrb SUBVID0_reg_5 ( .CK(PCICLK), .D(SUBVID02822_5), .R(HRST_), .QN(
        n6778) );
    zdffrb DEBUGC_reg_5 ( .CK(PCICLK), .D(DEBUGC3325_5), .R(HRST_), .QN(n6961)
         );
    zdffrb SUBSID0_reg_0 ( .CK(PCICLK), .D(SUBSID02898_0), .R(HRST_), .Q(
        SUBSID0_0), .QN(n6800) );
    zdffsb DEBUG8_reg_7 ( .CK(PCICLK), .D(DEBUG83126_7), .S(HRST_), .Q(
        DISCHKEOPERR), .QN(n6983) );
    zdffrb DEBUGB_reg_5 ( .CK(PCICLK), .D(DEBUGB3287_5), .R(HRST_), .Q(
        SLEEPTIME_SEL), .QN(n6969) );
    zdffrb SUBVID1_reg_5 ( .CK(PCICLK), .D(SUBVID12860_5), .R(HRST_), .QN(
        n6770) );
    zdffrb RxData_F_reg ( .CK(PCICLK), .D(RxData_F4946), .R(HRST_), .Q(
        RxData_F), .QN(n6805) );
    zdffqrb BIST_PATTERN_reg4_26 ( .CK(PCICLK), .D(n_11546), .R(HRST_), .Q(
        BIST_PATTERN[26]) );
    zivb U2147 ( .A(BIST_PATTERN[26]), .Y(n6710) );
    zdffrb SLQUEUE_ADDR_reg4_26 ( .CK(PCICLK), .D(n_6728), .R(HRST_), .Q(
        SLQUEUEADDR[26]), .QN(n6653) );
    zdffrb LAT_TM_reg_3 ( .CK(PCICLK), .D(LAT_TM2299_3), .R(HRST_), .QN(n6892)
         );
    zdffrb DEBUGD_reg_4 ( .CK(PCICLK), .D(DEBUGD3363_4), .R(HRST_), .QN(n6954)
         );
    zdffqrb Disconnect_H_reg ( .CK(PCICLK), .D(Disconnect_H5104), .R(HRST_), 
        .Q(Disconnect_H) );
    zdffrb PHYOPTEF_reg_1 ( .CK(PCICLK), .D(PHYOPTEF3629_1), .R(HRST_), .Q(
        CTRL_F[1]), .QN(n6842) );
    zdffrb TMOUT_PARM_reg_2 ( .CK(PCICLK), .D(TMOUT_PARM4236_2), .R(CMDRST_), 
        .Q(TMOUT_PARM[2]), .QN(n6738) );
    zdffqrb BIST_PATTERN_reg3_22 ( .CK(PCICLK), .D(n_10878), .R(HRST_), .Q(
        BIST_PATTERN[22]) );
    zivb U2148 ( .A(BIST_PATTERN[22]), .Y(n6716) );
    zdffrb SLQUEUE_ADDR_reg3_22 ( .CK(PCICLK), .D(n_6190), .R(HRST_), .Q(
        SLQUEUEADDR[22]), .QN(n6675) );
    zdffrb PHYOPT2_reg_6 ( .CK(PCICLK), .D(PHYOPT23515_6), .R(HRST_), .Q(
        SetPowner_Dis), .QN(n6862) );
    zdffqrb BIST_PATTERN_reg_0 ( .CK(PCICLK), .D(n_9570), .R(HRST_), .Q(
        BIST_PATTERN[0]) );
    zdffsb PHYOPT4_reg_7 ( .CK(PCICLK), .D(PHYOPT43591_7), .S(HRST_), .Q(
        CTRL_A[3]), .QN(n6845) );
    zdffrb IOBA10_reg ( .CK(PCICLK), .D(IOBA102699), .R(HRST_), .Q(IOBA10), 
        .QN(n6920) );
    zdffqrb BIST_PATTERN_reg2_14 ( .CK(PCICLK), .D(n_10218), .R(HRST_), .Q(
        BIST_PATTERN[14]) );
    zdffrb SUBVID0_reg_7 ( .CK(PCICLK), .D(SUBVID02822_7), .R(HRST_), .QN(
        n6776) );
    zdffrb DEBUGC_reg_7 ( .CK(PCICLK), .D(DEBUGC3325_7), .R(HRST_), .QN(n6959)
         );
    zdffrb SLQUEUE_ADDR_reg_2 ( .CK(PCICLK), .D(n_5142), .R(HRST_), .Q(
        SLQUEUEADDR[2]), .QN(n6693) );
    zdffrb SLQUEUE_ADDR_reg2_14 ( .CK(PCICLK), .D(n_5660), .R(HRST_), .Q(
        SLQUEUEADDR[14]), .QN(n6690) );
    zdffrb Squelch_E_reg ( .CK(PCICLK), .D(Squelch_E4855), .R(HRST_), .Q(
        Squelch_E), .QN(n6760) );
    zdffrb IOBA15_reg ( .CK(PCICLK), .D(IOBA152729), .R(HRST_), .Q(IOBA15), 
        .QN(n6915) );
    zdffrb SUBSID1_reg_2 ( .CK(PCICLK), .D(SUBSID12936_2), .R(HRST_), .QN(
        n6790) );
    zdffrb IOBA28_reg ( .CK(PCICLK), .D(IOBA282413), .R(HRST_), .Q(IOBA28), 
        .QN(n6902) );
    zdffrb PHYOPT3_reg_4 ( .CK(PCICLK), .D(PHYOPT33553_4), .R(HRST_), .Q(
        CTRL_C[0]), .QN(n6856) );
    zdffrb PHYOPT1_reg_0 ( .CK(PCICLK), .D(PHYOPT13477_0), .R(HRST_), .Q(CP0), 
        .QN(n6876) );
    zdffrb PHYOPTGH_reg_2 ( .CK(PCICLK), .D(PHYOPTGH3667_2), .R(HRST_), .Q(
        CTRL_H[2]), .QN(n6833) );
    zdffqrb SRAM_ADDR_IN_reg_5 ( .CK(PCICLK), .D(n_8044), .R(HRST_), .Q(
        SRAM_ADDR_IN_5) );
    zdffsb DEBUG2_reg_0 ( .CK(PCICLK), .D(DEBUG23050_0), .S(HRST_), .Q(
        OCUPY_SEL[0]), .QN(n7006) );
    zdffqrb RxData_C_reg ( .CK(PCICLK), .D(RxData_C4691), .R(HRST_), .Q(
        RxData_C) );
    zdffrb INTR_DIS_reg ( .CK(PCICLK), .D(INTR_DIS2113), .R(HRST_), .Q(
        INTR_DIS), .QN(n6921) );
    zdffrb PHYOPT4_reg_5 ( .CK(PCICLK), .D(PHYOPT43591_5), .R(HRST_), .Q(
        CTRL_A[1]), .QN(n6847) );
    zdffrb Disconnect_C_reg ( .CK(PCICLK), .D(Disconnect_C4679), .R(HRST_), 
        .Q(Disconnect_C), .QN(n6928) );
    zdffrb PHYOPT2_reg_4 ( .CK(PCICLK), .D(PHYOPT23515_4), .R(HRST_), .Q(
        RDOUT_Enb), .QN(n6864) );
    zdffrb SLQUEUE_ADDR_reg2_8 ( .CK(PCICLK), .D(n_5672), .R(HRST_), .Q(
        SLQUEUEADDR[8]), .QN(n6678) );
    zdffqrb BIST_PATTERN_reg_2 ( .CK(PCICLK), .D(n_9566), .R(HRST_), .Q(
        BIST_PATTERN[2]) );
    zdffrb RxDataDly_reg_1 ( .CK(PCICLK), .D(RxDataDly3781_1), .R(HRST_), .Q(
        RxDataDly[1]), .QN(n6811) );
    zdffrb SLQUEUE_ADDR_reg3_20 ( .CK(PCICLK), .D(n_6194), .R(HRST_), .Q(
        SLQUEUEADDR[20]), .QN(n6671) );
    zdffqrb BIST_PATTERN_reg3_20 ( .CK(PCICLK), .D(n_10882), .R(HRST_), .Q(
        BIST_PATTERN[20]) );
    zivb U2149 ( .A(BIST_PATTERN[20]), .Y(n6714) );
    zdffsb PHYOPTEF_reg_3 ( .CK(PCICLK), .D(PHYOPTEF3629_3), .S(HRST_), .Q(
        CTRL_F[3]), .QN(n6840) );
    zdffrb TMOUT_PARM_reg_0 ( .CK(PCICLK), .D(TMOUT_PARM4236_0), .R(CMDRST_), 
        .Q(TMOUT_PARM[0]), .QN(n6740) );
    zdffrb SLQUEUE_ADDR_reg4_24 ( .CK(PCICLK), .D(n_6732), .R(HRST_), .Q(
        SLQUEUEADDR[24]), .QN(n6649) );
    zdffrb CACHLN5_reg ( .CK(PCICLK), .D(CACHLN52194), .R(HRST_), .Q(CACHLN5), 
        .QN(n7029) );
    zdffsb LAT_TM_reg_1 ( .CK(PCICLK), .D(LAT_TM2299_1), .S(HRST_), .QN(n6894)
         );
    zdffrb DEBUGD_reg_6 ( .CK(PCICLK), .D(DEBUGD3363_6), .R(HRST_), .Q(
        DEBUGD_6), .QN(n6952) );
    zdffrb IOBA26_reg ( .CK(PCICLK), .D(IOBA262401), .R(HRST_), .Q(IOBA26), 
        .QN(n6904) );
    zdffqrb BIST_PATTERN_reg4_24 ( .CK(PCICLK), .D(n_11550), .R(HRST_), .Q(
        BIST_PATTERN[24]) );
    zdffrb DEBUGB_reg_7 ( .CK(PCICLK), .D(DEBUGB3287_7), .R(HRST_), .QN(n6967)
         );
    zdffrb SUBVID1_reg_7 ( .CK(PCICLK), .D(SUBVID12860_7), .R(HRST_), .QN(
        n6768) );
    zdffrb PHYMON_EN_E_reg ( .CK(PCICLK), .D(PHYMON_EN_E4386), .R(HRST_), .Q(
        PHYMON_EN_E), .QN(n6749) );
    zdffqrb SLAVEMODE_reg ( .CK(PCICLK_FREE), .D(SLAVEMODE4162), .R(CMDRST_), 
        .Q(SLAVEMODE) );
    zivb U2150 ( .A(SLAVEMODE), .Y(n6802) );
    zdffsb DEBUG8_reg_5 ( .CK(PCICLK), .D(DEBUG83126_5), .S(HRST_), .Q(
        DIS_BURST), .QN(n6985) );
    zdffsb SUBSID0_reg_2 ( .CK(PCICLK), .D(SUBSID02898_2), .S(HRST_), .Q(
        SUBSID0_2), .QN(n6798) );
    zdffqrb TERMON_A_reg ( .CK(PCICLK), .D(TERMON_A4503), .R(HRST_), .Q(
        TERMON_A) );
    zdffqrb TERMON_E_reg ( .CK(PCICLK), .D(TERMON_E4843), .R(HRST_), .Q(
        TERMON_E) );
    zdffsb DEBUG8_reg_2 ( .CK(PCICLK), .D(DEBUG83126_2), .S(HRST_), .Q(
        EN_UTM_RESET), .QN(n6988) );
    zdffrb SUBSID0_reg_5 ( .CK(PCICLK), .D(SUBSID02898_5), .R(HRST_), .Q(
        SUBSID0_5), .QN(n6795) );
    zdffsb DEBUGD_reg_1 ( .CK(PCICLK), .D(DEBUGD3363_1), .S(HRST_), .Q(
        EN_UTM_SPDUP), .QN(n6957) );
    zdffrb LAT_TM_reg_6 ( .CK(PCICLK), .D(LAT_TM2299_6), .R(HRST_), .Q(
        LAT_TM_6), .QN(n6889) );
    zdffrb IOBA22_reg ( .CK(PCICLK), .D(IOBA222574), .R(HRST_), .Q(IOBA22), 
        .QN(n6908) );
    zdffrb PHYMON_EN_A_reg ( .CK(PCICLK), .D(PHYMON_EN_A4362), .R(HRST_), .Q(
        PHYMON_EN_A), .QN(n6756) );
    zdffsb SUBVID1_reg_0 ( .CK(PCICLK), .D(SUBVID12860_0), .S(HRST_), .Q(
        SUBVID1_0), .QN(n6775) );
    zdffsb DEBUGB_reg_0 ( .CK(PCICLK), .D(DEBUGB3287_0), .S(HRST_), .Q(
        TURN_PARM[0]), .QN(n6974) );
    zdffrb CACHLN1_reg ( .CK(PCICLK), .D(CACHLN12170), .R(HRST_), .Q(CACHLN1), 
        .QN(n7042) );
    zdffqrb BACK_EN_reg ( .CK(PCICLK), .D(BACK_EN5715), .R(HRST_), .Q(BACK_EN)
         );
    zivb U2151 ( .A(BACK_EN), .Y(n7025) );
    zdffrb PHYOPTEF_reg_4 ( .CK(PCICLK), .D(PHYOPTEF3629_4), .R(HRST_), .Q(
        CTRL_E[0]), .QN(n6839) );
    zdffrb TMOUT_PARM_reg_7 ( .CK(PCICLK), .D(TMOUT_PARM4236_7), .R(CMDRST_), 
        .Q(TMOUT_PARM[7]), .QN(n6733) );
    zdffrb SRAM_WR_reg ( .CK(PCICLK), .D(SRAM_WR5337), .R(HRST_), .Q(SRAM_WR), 
        .QN(n6616) );
    zdffrb PHYOPT4_reg_2 ( .CK(PCICLK), .D(PHYOPT43591_2), .R(HRST_), .Q(
        CTRL_B[2]), .QN(n6850) );
    zdffrb Disconnect_G_reg ( .CK(PCICLK), .D(Disconnect_G5019), .R(HRST_), 
        .Q(Disconnect_G), .QN(n6925) );
    zdffqrb BIST_PATTERN_reg_5 ( .CK(PCICLK), .D(n_9560), .R(HRST_), .Q(
        BIST_PATTERN[5]) );
    zivb U2152 ( .A(BIST_PATTERN[5]), .Y(n6625) );
    zdffsb PHYOPT2_reg_3 ( .CK(PCICLK), .D(PHYOPT23515_3), .S(HRST_), .Q(
        FastLock), .QN(n6865) );
    zdffrb PHYOPTGH_reg_5 ( .CK(PCICLK), .D(PHYOPTGH3667_5), .R(HRST_), .Q(
        CTRL_G[1]), .QN(n6830) );
    zdffqrb SRAM_ADDR_IN_reg_2 ( .CK(PCICLK), .D(n_8050), .R(HRST_), .Q(
        SRAM_ADDR_IN_2) );
    zdffrb RxData_G_reg ( .CK(PCICLK), .D(RxData_G5031), .R(HRST_), .Q(
        RxData_G), .QN(n6804) );
    zdffrb PHYOPT1_reg_7 ( .CK(PCICLK), .D(PHYOPT13477_7), .R(HRST_), .Q(
        tst_buferr), .QN(n6869) );
    zdffrb DEBUG2_reg_7 ( .CK(PCICLK), .D(DEBUG23050_7), .R(HRST_), .Q(SELEOF), 
        .QN(n7000) );
    zdffsb PHYOPT3_reg_3 ( .CK(PCICLK), .D(PHYOPT33553_3), .S(HRST_), .Q(
        CTRL_D[3]), .QN(n6857) );
    zdffrb IOBA11_reg ( .CK(PCICLK), .D(IOBA112705), .R(HRST_), .Q(IOBA11), 
        .QN(n6919) );
    zdffrb DEBUG9_reg_2 ( .CK(PCICLK), .D(n_2804), .R(HRST_), .QN(n6705) );
    zdffqrb BIST_PATTERN_reg4_31 ( .CK(PCICLK), .D(n_11536), .R(HRST_), .Q(
        BIST_PATTERN[31]) );
    zdffsb SUBSID1_reg_5 ( .CK(PCICLK), .D(SUBSID12936_5), .S(HRST_), .Q(
        SUBSID1_5), .QN(n6787) );
    zdffqrb Squelch_A_reg ( .CK(PCICLK), .D(Squelch_A4515), .R(HRST_), .Q(
        Squelch_A) );
    zdffrb SLQUEUE_ADDR_reg4_31 ( .CK(PCICLK), .D(n_6718), .R(HRST_), .Q(
        SLQUEUEADDR[31]), .QN(n6660) );
    zdffrb BMASTREN_reg ( .CK(PCICLK), .D(BMASTREN2046), .R(HRST_), .Q(
        BMASTREN), .QN(n7041) );
    zdffrb SLQUEUE_ADDR_reg2_13 ( .CK(PCICLK), .D(n_5662), .R(HRST_), .Q(
        SLQUEUEADDR[13]), .QN(n6688) );
    zdffrb SLQUEUE_ADDR_reg_5 ( .CK(PCICLK), .D(n_5136), .R(HRST_), .Q(
        SLQUEUEADDR[5]), .QN(n6696) );
    zdffrb SUBVID0_reg_0 ( .CK(PCICLK), .D(SUBVID02822_0), .R(HRST_), .Q(
        SUBVID0_0), .QN(n6783) );
    zdffrb DEBUGC_reg_0 ( .CK(PCICLK), .D(DEBUGC3325_0), .R(HRST_), .Q(SQSET
        [0]), .QN(n6966) );
    zdffqrb BIST_PATTERN_reg2_13 ( .CK(PCICLK), .D(n_10220), .R(HRST_), .Q(
        BIST_PATTERN[13]) );
    zivb U2153 ( .A(BIST_PATTERN[13]), .Y(n6720) );
    zdffsb PHYOPT4_reg_3 ( .CK(PCICLK), .D(PHYOPT43591_3), .S(HRST_), .Q(
        CTRL_B[3]), .QN(n6849) );
    zdffqrb BIST_PATTERN_reg_4 ( .CK(PCICLK), .D(n_9562), .R(HRST_), .Q(
        BIST_PATTERN[4]) );
    zivb U2154 ( .A(BIST_PATTERN[4]), .Y(n6623) );
    zdffrb IOBA19_reg ( .CK(PCICLK), .D(IOBA192556), .R(HRST_), .Q(IOBA19), 
        .QN(n6911) );
    zdffrb PHYOPT2_reg_2 ( .CK(PCICLK), .D(PHYOPT23515_2), .R(HRST_), .Q(
        LBack_Enb), .QN(n6866) );
    zdffrb Disconnect_A_reg ( .CK(PCICLK), .D(Disconnect_A4509), .R(HRST_), 
        .Q(Disconnect_A), .QN(n6930) );
    zdffrb PHYOPTEF_reg_5 ( .CK(PCICLK), .D(PHYOPTEF3629_5), .R(HRST_), .Q(
        CTRL_E[1]), .QN(n6838) );
    zdffsb TMOUT_PARM_reg_6 ( .CK(PCICLK), .D(TMOUT_PARM4236_6), .S(CMDRST_), 
        .Q(TMOUT_PARM[6]), .QN(n6734) );
    zdffrb TERMON_C_reg ( .CK(PCICLK), .D(TERMON_C4673), .R(HRST_), .Q(
        TERMON_C), .QN(n6753) );
    zdffrb LAT_TM_reg_7 ( .CK(PCICLK), .D(LAT_TM2299_7), .R(HRST_), .QN(n6888)
         );
    zdffsb DEBUGD_reg_0 ( .CK(PCICLK), .D(DEBUGD3363_0), .S(HRST_), .Q(
        EN_DBG_PORT), .QN(n6958) );
    zdffrb SUBVID1_reg_1 ( .CK(PCICLK), .D(SUBVID12860_1), .R(HRST_), .QN(
        n6774) );
    zdffrb DEBUGB_reg_1 ( .CK(PCICLK), .D(DEBUGB3287_1), .R(HRST_), .Q(
        TURN_PARM[1]), .QN(n6973) );
    zdffrb PHYMON_EN_G_reg ( .CK(PCICLK), .D(PHYMON_EN_G4398), .R(HRST_), .Q(
        PHYMON_EN_G), .QN(n6747) );
    zdffrb DEBUG8_reg_3 ( .CK(PCICLK), .D(DEBUG83126_3), .R(HRST_), .Q(
        DISPSTUFF), .QN(n6987) );
    zdffrb IOBA24_reg ( .CK(PCICLK), .D(IOBA242389), .R(HRST_), .Q(IOBA24), 
        .QN(n6906) );
    zdffrb SUBSID0_reg_4 ( .CK(PCICLK), .D(SUBSID02898_4), .R(HRST_), .Q(
        SUBSID0_4), .QN(n6796) );
    zdffrb CACHLN7_reg ( .CK(PCICLK), .D(CACHLN72206), .R(HRST_), .Q(CACHLN7), 
        .QN(n7027) );
    zdffrb IOBA8_reg ( .CK(PCICLK), .D(IOBA82687), .R(HRST_), .Q(IOBA8), .QN(
        n6898) );
    zdffrb IOBA30_reg ( .CK(PCICLK), .D(IOBA302425), .R(HRST_), .Q(IOBA30), 
        .QN(n6900) );
    zdffrb IOBA17_reg ( .CK(PCICLK), .D(IOBA172544), .R(HRST_), .Q(IOBA17), 
        .QN(n6913) );
    zdffrb SLQUEUE_ADDR_reg2_12 ( .CK(PCICLK), .D(n_5664), .R(HRST_), .Q(
        SLQUEUEADDR[12]), .QN(n6686) );
    zdffrb SLQUEUE_ADDR_reg_4 ( .CK(PCICLK), .D(n_5138), .R(HRST_), .Q(
        SLQUEUEADDR[4]), .QN(n6695) );
    zdffsb DEBUGC_reg_1 ( .CK(PCICLK), .D(DEBUGC3325_1), .S(HRST_), .Q(SQSET
        [1]), .QN(n6965) );
    zdffrb Squelch_G_reg ( .CK(PCICLK), .D(Squelch_G5025), .R(HRST_), .Q(
        Squelch_G), .QN(n6758) );
    zdffqrb BIST_PATTERN_reg2_12 ( .CK(PCICLK), .D(n_10222), .R(HRST_), .Q(
        BIST_PATTERN[12]) );
    zivb U2155 ( .A(BIST_PATTERN[12]), .Y(n6719) );
    zdffrb DEBUG9_reg_3 ( .CK(PCICLK), .D(n_2802), .R(HRST_), .QN(n6706) );
    zdffqrb BIST_PATTERN_reg4_30 ( .CK(PCICLK), .D(n_11538), .R(HRST_), .Q(
        BIST_PATTERN[30]) );
    zdffsb SUBSID1_reg_4 ( .CK(PCICLK), .D(SUBSID12936_4), .S(HRST_), .Q(
        SUBSID1_4), .QN(n6788) );
    zdffrb SLQUEUE_ADDR_reg4_30 ( .CK(PCICLK), .D(n_6720), .R(HRST_), .Q(
        SLQUEUEADDR[30]), .QN(n6658) );
    zdffrb RxData_A_reg ( .CK(PCICLK), .D(RxData_A4521), .R(HRST_), .Q(
        RxData_A), .QN(n6809) );
    zdffrb PHYOPT3_reg_2 ( .CK(PCICLK), .D(PHYOPT33553_2), .R(HRST_), .Q(
        CTRL_D[2]), .QN(n6858) );
    zdffrb PHYOPTGH_reg_4 ( .CK(PCICLK), .D(PHYOPTGH3667_4), .R(HRST_), .Q(
        CTRL_G[0]), .QN(n6831) );
    zdffqrb SRAM_ADDR_IN_reg_3 ( .CK(PCICLK), .D(n_8048), .R(HRST_), .Q(
        SRAM_ADDR_IN_3) );
    zdffrb PHYOPT1_reg_6 ( .CK(PCICLK), .D(PHYOPT13477_6), .R(HRST_), .Q(
        FAST_RST), .QN(n6870) );
    zdffrb DEBUG2_reg_6 ( .CK(PCICLK), .D(DEBUG23050_6), .R(HRST_), .Q(
        ENTXDLY_3), .QN(n7001) );
    zdffrb PHYOPT1_reg_1 ( .CK(PCICLK), .D(PHYOPT13477_1), .R(HRST_), .Q(CP1), 
        .QN(n6875) );
    zdffsb PHYOPTGH_reg_3 ( .CK(PCICLK), .D(PHYOPTGH3667_3), .S(HRST_), .Q(
        CTRL_H[3]), .QN(n6832) );
    zdffqrb SRAM_ADDR_IN_reg_4 ( .CK(PCICLK), .D(n_8046), .R(HRST_), .Q(
        SRAM_ADDR_IN_4) );
    zdffrb MMSPACE_reg ( .CK(PCICLK), .D(MMSPACE2040), .R(HRST_), .Q(MMSPACE), 
        .QN(n6885) );
    zdffsb DEBUG2_reg_1 ( .CK(PCICLK), .D(DEBUG23050_1), .S(HRST_), .Q(
        OCUPY_SEL[1]), .QN(n7005) );
    zdffrb MWRMEN_reg ( .CK(PCICLK), .D(MWRMEN2052), .R(HRST_), .Q(MWRMEN), 
        .QN(n6884) );
    zdffrb PHYOPT3_reg_5 ( .CK(PCICLK), .D(PHYOPT33553_5), .R(HRST_), .Q(
        CTRL_C[1]), .QN(n6855) );
    zdffrb RxData_E_reg ( .CK(PCICLK), .D(RxData_E4861), .R(HRST_), .Q(
        RxData_E), .QN(n6806) );
    zdffsb CLKOFF_EN_reg ( .CK(PCICLK_FREE), .D(CLKOFF_EN3164), .S(HRST_), .Q(
        CLKOFF_EN), .QN(n7020) );
    zdffrb DEBUG9_reg_4 ( .CK(PCICLK), .D(n_2800), .R(HRST_), .Q(DISPDRCV), 
        .QN(n6707) );
    zdffrb SUBSID1_reg_3 ( .CK(PCICLK), .D(SUBSID12936_3), .R(HRST_), .QN(
        n6789) );
    zdffrb Squelch_C_reg ( .CK(PCICLK), .D(Squelch_C4685), .R(HRST_), .Q(
        Squelch_C), .QN(n6762) );
    zdffqrb SLAVE_ACT_T_reg ( .CK(PCICLK_FREE), .D(SLAVE_ACT), .R(CMDRST_), 
        .Q(SLAVE_ACT_T) );
    zdffqrb BIST_PATTERN_reg2_15 ( .CK(PCICLK), .D(n_10216), .R(HRST_), .Q(
        BIST_PATTERN[15]) );
    zdffrb SUBVID0_reg_6 ( .CK(PCICLK), .D(SUBVID02822_6), .R(HRST_), .QN(
        n6777) );
    zdffrb DEBUGC_reg_6 ( .CK(PCICLK), .D(DEBUGC3325_6), .R(HRST_), .QN(n6960)
         );
    zdffrb IOBA13_reg ( .CK(PCICLK), .D(IOBA132717), .R(HRST_), .Q(IOBA13), 
        .QN(n6917) );
    zdffrb SLQUEUE_ADDR_reg_3 ( .CK(PCICLK), .D(n_5140), .R(HRST_), .Q(
        SLQUEUEADDR[3]), .QN(n6694) );
    zdffrb SLQUEUE_ADDR_reg2_15 ( .CK(PCICLK), .D(n_5658), .R(HRST_), .Q(
        SLQUEUEADDR[15]), .QN(n6692) );
    zdffrb CACHLN3_reg ( .CK(PCICLK), .D(CACHLN32182), .R(HRST_), .Q(CACHLN3), 
        .QN(n7033) );
    zdffsb DEBUG8_reg_4 ( .CK(PCICLK), .D(DEBUG83126_4), .S(HRST_), .Q(
        EN_REF_RVLD), .QN(n6986) );
    zdffrb IOBA20_reg ( .CK(PCICLK), .D(IOBA202562), .R(HRST_), .Q(IOBA20), 
        .QN(n6910) );
    zdffrb PHYMON_EN_C_reg ( .CK(PCICLK), .D(PHYMON_EN_C4374), .R(HRST_), .Q(
        PHYMON_EN_C), .QN(n6752) );
    zdffrb SUBSID0_reg_3 ( .CK(PCICLK), .D(SUBSID02898_3), .R(HRST_), .Q(
        SUBSID0_3), .QN(n6797) );
    zdffrb SLQUEUE_ADDR_reg4_25 ( .CK(PCICLK), .D(n_6730), .R(HRST_), .Q(
        SLQUEUEADDR[25]), .QN(n6651) );
    zdffrb DEBUGD_reg_7 ( .CK(PCICLK), .D(DEBUGD3363_7), .R(HRST_), .QN(n6951)
         );
    zdffrb LAT_TM_reg_0 ( .CK(PCICLK), .D(LAT_TM2299_0), .R(HRST_), .Q(
        LAT_TM_0), .QN(n6895) );
    zdffqrb BIST_PATTERN_reg4_25 ( .CK(PCICLK), .D(n_11548), .R(HRST_), .Q(
        BIST_PATTERN[25]) );
    zdffrb SUBVID1_reg_6 ( .CK(PCICLK), .D(SUBVID12860_6), .R(HRST_), .QN(
        n6769) );
    zdffrb DEBUGB_reg_6 ( .CK(PCICLK), .D(DEBUGB3287_6), .R(HRST_), .Q(
        DIS_NARROW_SOF), .QN(n6968) );
    zdffrb SWDBG_reg ( .CK(PCICLK), .D(SWDBG4088), .R(CMDRST_), .Q(SWDBG), 
        .QN(n6430) );
    zdffqrb TERMON_G_reg ( .CK(PCICLK), .D(TERMON_G5013), .R(HRST_), .Q(
        TERMON_G) );
    zdffrb SLQUEUE_ADDR_reg3_21 ( .CK(PCICLK), .D(n_6192), .R(HRST_), .Q(
        SLQUEUEADDR[21]), .QN(n6673) );
    zdffqrb BIST_PATTERN_reg3_21 ( .CK(PCICLK), .D(n_10880), .R(HRST_), .Q(
        BIST_PATTERN[21]) );
    zivb U2156 ( .A(BIST_PATTERN[21]), .Y(n6715) );
    zdffrb FastStart_reg ( .CK(PCICLK), .D(FastStart3819), .R(HRST_), .Q(
        FastStart), .QN(n6923) );
    zdffrb Disconnect_E_reg ( .CK(PCICLK), .D(Disconnect_E4849), .R(HRST_), 
        .Q(Disconnect_E), .QN(n6926) );
    zdffrb PHYOPTEF_reg_2 ( .CK(PCICLK), .D(PHYOPTEF3629_2), .R(HRST_), .Q(
        CTRL_F[2]), .QN(n6841) );
    zdffrb TMOUT_PARM_reg_1 ( .CK(PCICLK), .D(TMOUT_PARM4236_1), .R(CMDRST_), 
        .Q(TMOUT_PARM[1]), .QN(n6739) );
    zdffrb PHYOPT4_reg_4 ( .CK(PCICLK), .D(PHYOPT43591_4), .R(HRST_), .Q(
        CTRL_A[0]), .QN(n6848) );
    zdffrb SLQUEUE_ADDR_reg2_9 ( .CK(PCICLK), .D(n_5670), .R(HRST_), .Q(
        SLQUEUEADDR[9]), .QN(n6680) );
    zdffrb PHYOPT2_reg_5 ( .CK(PCICLK), .D(PHYOPT23515_5), .R(HRST_), .Q(
        autochk), .QN(n6863) );
    zdffsb RxDataDly_reg_0 ( .CK(PCICLK), .D(RxDataDly3781_0), .S(HRST_), .Q(
        RxDataDly[0]), .QN(n6812) );
    zdffqrb BIST_PATTERN_reg_3 ( .CK(PCICLK), .D(n_9564), .R(HRST_), .Q(
        BIST_PATTERN[3]) );
    zivb U2157 ( .A(BIST_PATTERN[3]), .Y(n6621) );
    znr2d U2158 ( .A(n6632), .B(n7140), .Y(n6337) );
    znr2d U2159 ( .A(n6661), .B(n6934), .Y(n6338) );
    znr2d U2160 ( .A(n6645), .B(n6765), .Y(n6339) );
    znr2d U2161 ( .A(n6661), .B(n7129), .Y(n6340) );
    znr2d U2162 ( .A(n7135), .B(n6661), .Y(n6342) );
    znr2b U2163 ( .A(n6661), .B(n7138), .Y(n6343) );
    znr2d U2164 ( .A(n6646), .B(n6991), .Y(n6344) );
    znr2b U2165 ( .A(n6661), .B(n6827), .Y(n6345) );
    znr2b U2166 ( .A(n6765), .B(n6878), .Y(n6346) );
    znr2d U2167 ( .A(n6632), .B(n7137), .Y(n6347) );
    znr2d U2168 ( .A(n7134), .B(n6632), .Y(n6348) );
    znr2b U2169 ( .A(n6632), .B(n6815), .Y(n6349) );
    znr2d U2170 ( .A(n6646), .B(n7131), .Y(n6350) );
    znr2d U2171 ( .A(n6646), .B(n7139), .Y(n6351) );
    znr2b U2172 ( .A(n6661), .B(n6702), .Y(n6352) );
    znr2d U2173 ( .A(n6614), .B(n6646), .Y(n6353) );
    znr2b U2174 ( .A(n6700), .B(n6765), .Y(n6354) );
    znr2b U2175 ( .A(n7140), .B(n6661), .Y(n6355) );
    znr2b U2176 ( .A(n6585), .B(n6764), .Y(n6356) );
    znr2b U2177 ( .A(n6633), .B(n6645), .Y(n6357) );
    znr2b U2178 ( .A(n6633), .B(n6700), .Y(n6358) );
    znr2b U2179 ( .A(n6646), .B(n6844), .Y(n6359) );
    znr2b U2180 ( .A(n6631), .B(n6878), .Y(n6360) );
    znr2d U2181 ( .A(n6729), .B(n6766), .Y(n6361) );
    znr2b U2182 ( .A(n6611), .B(n6824), .Y(n6362) );
    znr3b U2183 ( .A(n6701), .B(n6958), .C(n6824), .Y(n6363) );
    znr2b U2184 ( .A(n7022), .B(n7023), .Y(n6364) );
    znr2b U2185 ( .A(n7031), .B(n7032), .Y(n6365) );
    znr2b U2186 ( .A(n6342), .B(n6615), .Y(n6366) );
    znr2b U2187 ( .A(n6342), .B(SRAM_LAT_RDATA), .Y(n6367) );
    znr2b U2188 ( .A(n6348), .B(n6615), .Y(n6368) );
    znr2b U2189 ( .A(n6348), .B(SRAM_LAT_RDATA), .Y(n6369) );
    znr2b U2190 ( .A(n6353), .B(n6615), .Y(n6370) );
    znr2b U2191 ( .A(n6436), .B(n6615), .Y(n6371) );
    znr2b U2192 ( .A(SRAM_LAT_RDATA), .B(n6353), .Y(n6372) );
    znr2d U2193 ( .A(SRAM_LAT_RDATA), .B(n6436), .Y(n6373) );
    znr2b U2194 ( .A(n7025), .B(n7026), .Y(n6374) );
    znr3d U2195 ( .A(n6767), .B(n6766), .C(n6765), .Y(n6375) );
    znr3d U2196 ( .A(n6767), .B(n6766), .C(n6730), .Y(n6376) );
    znr3d U2197 ( .A(n6784), .B(n6767), .C(n6646), .Y(n6377) );
    znr3d U2198 ( .A(n7136), .B(n6767), .C(n6661), .Y(n6378) );
    znr2b U2199 ( .A(n6635), .B(n6646), .Y(n6379) );
    znr2b U2200 ( .A(n6632), .B(n6879), .Y(n6380) );
    znr2b U2201 ( .A(n6613), .B(n6879), .Y(n6381) );
    znr2d U2202 ( .A(n6633), .B(n6880), .Y(n6382) );
    znr2d U2203 ( .A(n6646), .B(n6881), .Y(n6383) );
    znr2d U2204 ( .A(n6661), .B(n6881), .Y(n6384) );
    ziv11b U2205 ( .A(n6146), .Y(n6385), .Z(n6386) );
    zivb U2206 ( .A(n6827), .Y(n6387) );
    zao22b U2207 ( .A(n7069), .B(TrkSpd[1]), .C(USBLEGSUP[3]), .D(n6422), .Y(
        n7088) );
    zao22b U2208 ( .A(n7069), .B(TERMON_G), .C(SUBSID1_0), .D(n6361), .Y(n6547
        ) );
    zao22b U2209 ( .A(LBack_Enb), .B(n7070), .C(CTRL_F[2]), .D(n7069), .Y(
        n6481) );
    zbfb U2210 ( .A(n6827), .Y(n6388) );
    zoai2x4b U2211 ( .A(n6388), .B(n6842), .C(n7139), .D(n6680), .E(n7127), 
        .F(n6930), .G(n6774), .H(n7136), .Y(n6476) );
    zoai2x4b U2212 ( .A(n6388), .B(n6839), .C(n7140), .D(n6686), .E(n6771), 
        .F(n6784), .G(n6755), .H(n6877), .Y(n6491) );
    zoai2x4b U2213 ( .A(n6388), .B(n6923), .C(n7129), .D(n7013), .E(n7139), 
        .F(n6698), .G(n7024), .H(n7027), .Y(n7077) );
    zoai2x4b U2214 ( .A(n6810), .B(n6827), .C(n7128), .D(n7014), .E(n6741), 
        .F(n6924), .G(n7139), .H(n6697), .Y(n6467) );
    zoai2x4b U2215 ( .A(n6811), .B(n6827), .C(n6741), .D(n6745), .E(n7129), 
        .F(n7015), .G(n6647), .H(n6696), .Y(n6463) );
    zoai2x4b U2216 ( .A(n7137), .B(n6863), .C(n6827), .D(n6838), .E(n6647), 
        .F(n6688), .G(n6770), .H(n7136), .Y(n6495) );
    zoai2x4b U2217 ( .A(n7137), .B(n6861), .C(n6827), .D(n6836), .E(n7140), 
        .F(n6692), .G(n6768), .H(n6784), .Y(n6506) );
    zoai2x4b U2218 ( .A(n6844), .B(n6865), .C(n6827), .D(n6840), .E(n7140), 
        .F(n6684), .G(n6809), .H(n7127), .Y(n6489) );
    zoai2x4b U2219 ( .A(n7138), .B(n6862), .C(n6827), .D(n6837), .E(n7139), 
        .F(n6690), .G(n6769), .H(n7136), .Y(n6499) );
    zoai2x4b U2220 ( .A(n6759), .B(n7127), .C(n6757), .D(n6827), .E(n7136), 
        .F(n6786), .G(n7132), .H(n6968), .Y(n6575) );
    zoai2x4b U2221 ( .A(n7138), .B(n6849), .C(n6804), .D(n6827), .E(n6784), 
        .F(n6789), .G(n6702), .H(n6971), .Y(n6559) );
    zoai2x4b U2222 ( .A(n7137), .B(n6850), .C(n6758), .D(n6827), .E(n7136), 
        .F(n6790), .G(n7133), .H(n6972), .Y(n6555) );
    zoai2x4b U2223 ( .A(n6805), .B(n6877), .C(n6803), .D(n6827), .E(n7136), 
        .F(n6785), .G(n7133), .H(n6967), .Y(n6579) );
    zoai2x4b U2224 ( .A(n6779), .B(n6784), .C(n6812), .D(n6827), .E(n7128), 
        .F(n7016), .G(n7140), .H(n6695), .Y(n6458) );
    zoai2x4b U2225 ( .A(n7129), .B(n6998), .C(n6934), .D(n6941), .E(n6844), 
        .F(n6851), .G(n6827), .H(n6925), .Y(n6552) );
    zivb U2226 ( .A(n6827), .Y(n7069) );
    zor2b U2227 ( .A(n6645), .B(n6729), .Y(n6827) );
    zivb U2228 ( .A(n6882), .Y(n6389) );
    zan2b U2229 ( .A(n6425), .B(n6420), .Y(PCI_R6FG) );
    zan2b U2230 ( .A(USBLEGCTLSTS[2]), .B(n6389), .Y(n6599) );
    zao2x4b U2231 ( .A(CACHLN6), .B(n7068), .C(USBLEGSUP[6]), .D(n6422), .E(
        USBLEGCTLSTS[6]), .F(n6389), .G(n6374), .H(REVID_BACK_6), .Y(n6466) );
    zao22b U2232 ( .A(USBLEGCTLSTS[0]), .B(n6389), .C(PWR_STATE0), .D(n6362), 
        .Y(n7111) );
    zao22b U2233 ( .A(USBLEGSUP[24]), .B(n6422), .C(USBLEGCTLSTS[24]), .D(
        n6425), .Y(n7092) );
    zao22b U2234 ( .A(USBLEGSUP[20]), .B(n6422), .C(USBLEGCTLSTS[20]), .D(
        n6389), .Y(n6528) );
    zao22b U2235 ( .A(USBLEGSUP[22]), .B(n6422), .C(USBLEGCTLSTS[22]), .D(
        n6389), .Y(n6538) );
    zivb U2236 ( .A(n6882), .Y(n6425) );
    zivb U2237 ( .A(n6882), .Y(n7125) );
    zivb U2238 ( .A(n6883), .Y(n6390) );
    zan2b U2239 ( .A(n6390), .B(n6417), .Y(PCI_R6AG) );
    zao2x4b U2240 ( .A(BIST_PATTERN[14]), .B(n7059), .C(IOBA14), .D(n6586), 
        .E(USBLEGSUP[14]), .F(n6422), .G(USBLEGCTLSTS[14]), .H(n6425), .Y(
        n6501) );
    zao22b U2241 ( .A(USBLEGSUP[18]), .B(n6390), .C(USBLEGCTLSTS[18]), .D(
        n6425), .Y(n6517) );
    zao22b U2242 ( .A(USBLEGSUP[23]), .B(n6390), .C(USBLEGCTLSTS[23]), .D(
        n6389), .Y(n7096) );
    zao22b U2243 ( .A(USBLEGSUP[8]), .B(n7124), .C(USBLEGCTLSTS[8]), .D(n6389), 
        .Y(n6474) );
    zao22b U2244 ( .A(USBLEGSUP[21]), .B(n7124), .C(USBLEGCTLSTS[21]), .D(
        n6425), .Y(n6533) );
    zao22b U2245 ( .A(n7069), .B(TrkSpd[0]), .C(USBLEGSUP[2]), .D(n7124), .Y(
        n6450) );
    zao22b U2246 ( .A(CACHLN5), .B(n7068), .C(USBLEGSUP[5]), .D(n6390), .Y(
        n7079) );
    zivb U2247 ( .A(n6883), .Y(n7124) );
    zivb U2248 ( .A(n6883), .Y(n6422) );
    zivb U2249 ( .A(n6741), .Y(n6391) );
    zao22b U2250 ( .A(CACHLN4), .B(n7068), .C(UTM_CHKERR), .D(n6391), .Y(n6457
        ) );
    zao22b U2251 ( .A(SL_ET_ERR), .B(n7062), .C(USBLEGSUP[19]), .D(n6390), .Y(
        n6525) );
    zao22b U2252 ( .A(PIDERR), .B(n7062), .C(USBLEGSUP[17]), .D(n7124), .Y(
        n7100) );
    zao22b U2253 ( .A(SL_ERROFFSET[4]), .B(n7062), .C(USBLEGSUP[28]), .D(n7124
        ), .Y(n6567) );
    zao22b U2254 ( .A(SL_ERROFFSET[1]), .B(n7062), .C(USBLEGSUP[25]), .D(n7124
        ), .Y(n7091) );
    zao22b U2255 ( .A(SL_ERROFFSET[6]), .B(n7062), .C(USBLEGSUP[30]), .D(n6390
        ), .Y(n7086) );
    zivb U2256 ( .A(n6741), .Y(n7062) );
    zor2b U2257 ( .A(n6631), .B(n6645), .Y(n6741) );
    zivb U2258 ( .A(n6826), .Y(n6392) );
    zan2b U2259 ( .A(n6392), .B(n6417), .Y(R62G) );
    zan2b U2260 ( .A(n6392), .B(n6420), .Y(R63G) );
    zao22b U2261 ( .A(FLADJ3), .B(n6416), .C(USBLEGCTLSTS[11]), .D(n6425), .Y(
        n6487) );
    zao22b U2262 ( .A(PORTWAKECAP0), .B(n6416), .C(USBLEGSUP[16]), .D(n6390), 
        .Y(n7103) );
    zao22b U2263 ( .A(IOBA8), .B(n6586), .C(FLADJ0), .D(n6416), .Y(n6472) );
    zan3b U2264 ( .A(PORTWAKECAP4), .B(ENUSB2), .C(n6416), .Y(n6598) );
    zan3b U2265 ( .A(PORTWAKECAP6), .B(ENUSB3), .C(n6416), .Y(n6596) );
    zan3b U2266 ( .A(ENUSB3), .B(PORTWAKECAP5), .C(n6416), .Y(n6597) );
    zan3b U2267 ( .A(PORTWAKECAP2), .B(ENUSB1), .C(n6416), .Y(n6600) );
    zan3b U2268 ( .A(PORTWAKECAP8), .B(ENUSB4), .C(n6416), .Y(n6595) );
    zao32b U2269 ( .A(ENUSB1), .B(PORTWAKECAP1), .C(n6416), .D(REVID1), .E(
        n7058), .Y(n7099) );
    zao21b U2270 ( .A(USBLEGCTLSTS[5]), .B(n6425), .C(n6416), .Y(n7078) );
    zor2b U2271 ( .A(n6631), .B(n6825), .Y(n6826) );
    zivb U2272 ( .A(n6826), .Y(n6416) );
    zivb U2273 ( .A(n7023), .Y(n6393) );
    zao22b U2274 ( .A(USBLEGCTLSTS[10]), .B(n6425), .C(n6393), .D(n7022), .Y(
        n6484) );
    zao2x4b U2275 ( .A(CTRL_H[2]), .B(n7069), .C(SUBSID0_2), .D(n6361), .E(
        MINGNT2), .F(n7084), .G(SL_DATA_PIDERR), .H(n7062), .Y(n6518) );
    zao2x4b U2276 ( .A(CTRL_G[1]), .B(n7069), .C(SUBSID0_5), .D(n6361), .E(
        MINGNT5), .F(n7084), .G(SL_ACK_ERR), .H(n7062), .Y(n6534) );
    zao2x4b U2277 ( .A(SLQUEUEADDR[24]), .B(n7065), .C(BIST_PATTERN[24]), .D(
        n7059), .E(MAXLAT0), .F(n7084), .G(SL_ERROFFSET[0]), .H(n7062), .Y(
        n6550) );
    zao2x4b U2278 ( .A(CTRL_H[0]), .B(n7069), .C(SUBSID0_0), .D(n6361), .E(
        MINGNT0), .F(n7084), .G(CRCERR), .H(n7062), .Y(n6511) );
    zao2x4b U2279 ( .A(CTRL_G[0]), .B(n7069), .C(SUBSID0_4), .D(n6361), .E(
        MINGNT4), .F(n7084), .G(SL_SE_ERR), .H(n7062), .Y(n6529) );
    zao2x4b U2280 ( .A(CTRL_G[2]), .B(n7069), .C(SUBSID0_6), .D(n6361), .E(
        MINGNT6), .F(n7084), .G(SL_PCIERR), .H(n7062), .Y(n6539) );
    zao2x4b U2281 ( .A(CTRL_H[3]), .B(n7069), .C(SUBSID0_3), .D(n6361), .E(
        UIRQACT), .F(n7083), .G(MINGNT3), .H(n7084), .Y(n6526) );
    zao2x4b U2282 ( .A(IOBA31), .B(n6586), .C(SLQUEUEADDR[31]), .D(n7065), .E(
        BIST_PATTERN[31]), .F(n7059), .G(MAXLAT7), .H(n7084), .Y(n6582) );
    zao2x4b U2283 ( .A(SLQUEUEADDR[25]), .B(n7065), .C(BIST_PATTERN[25]), .D(
        n7059), .E(DEVS0), .F(n7083), .G(MAXLAT1), .H(n7084), .Y(n6554) );
    zao2x4b U2284 ( .A(BIST_PATTERN[17]), .B(n7059), .C(CTRL_H[1]), .D(n7069), 
        .E(SUBSID0_1), .F(n6361), .G(MINGNT1), .H(n7084), .Y(n6515) );
    zao2x4b U2285 ( .A(IOBA30), .B(n6586), .C(SLQUEUEADDR[30]), .D(n7065), .E(
        BIST_PATTERN[30]), .F(n7059), .G(MAXLAT6), .H(n7084), .Y(n6578) );
    zao2x4b U2286 ( .A(IOBA28), .B(n6586), .C(SLQUEUEADDR[28]), .D(n7065), .E(
        BIST_PATTERN[28]), .F(n7059), .G(MAXLAT4), .H(n7084), .Y(n6568) );
    zao2x4b U2287 ( .A(MAXLAT2), .B(n7084), .C(SL_ERROFFSET[2]), .D(n7062), 
        .E(USBLEGSUP[26]), .F(n6422), .G(USBLEGCTLSTS[26]), .H(n6425), .Y(
        n6557) );
    zao2x4b U2288 ( .A(MAXLAT3), .B(n7084), .C(SL_ERROFFSET[3]), .D(n7062), 
        .E(USBLEGSUP[27]), .F(n6390), .G(USBLEGCTLSTS[27]), .H(n6389), .Y(
        n6561) );
    zor2b U2289 ( .A(n6729), .B(n6922), .Y(n7023) );
    zivb U2290 ( .A(n7023), .Y(n7084) );
    zbfd U2291 ( .A(n6146), .Y(SRAM_SEL[1]) );
    zbfd U2292 ( .A(n6146), .Y(n6395) );
    zdffqrb SRAM_SEL_reg_1 ( .CK(PCICLK), .D(SRAM_SEL5343_1), .R(HRST_), .Q(
        n6146) );
    zbfd U2293 ( .A(n6145), .Y(SRAM_SEL[0]) );
    zbfb U2294 ( .A(n6145), .Y(n6397) );
    zivb U2295 ( .A(n6145), .Y(n6801) );
    zdffqrb SRAM_SEL_reg_0 ( .CK(PCICLK), .D(SRAM_SEL5343_0), .R(HRST_), .Q(
        n6145) );
    zor2b U2296 ( .A(CBE0I_), .B(n6741), .Y(n6398) );
    znr2b U2297 ( .A(CBE0I_), .B(n6612), .Y(n6399) );
    zivb U2298 ( .A(n6399), .Y(n6613) );
    zivb U2299 ( .A(CFGW), .Y(n6612) );
    zdffsd SUBVID0_reg_1 ( .CK(PCICLK), .D(SUBVID02822_1), .S(HRST_), .Q(
        SUBVID0_1), .QN(n6782) );
    zan2d U2300 ( .A(n6419), .B(n6415), .Y(n6418) );
    zan2d U2301 ( .A(n7124), .B(n6420), .Y(PCI_R6BG) );
    zor4b U2302 ( .A(n6384), .B(n6424), .C(n6383), .D(n6382), .Y(PCI_RBAR) );
    zan2d U2303 ( .A(n6362), .B(n6426), .Y(R85G) );
    zan4b U2304 ( .A(n6429), .B(n6430), .C(n6431), .D(n6432), .Y(n6428) );
    zan2d U2305 ( .A(n6434), .B(n6435), .Y(BIST_ERROR4199) );
    zao222b U2306 ( .A(SRAM_RDATA_SEL_7), .B(n6371), .C(BIST_PATTERN[7]), .D(
        n6373), .E(AD7I), .F(n6436), .Y(n_9556) );
    zao222b U2307 ( .A(SRAM_RDATA_SEL_6), .B(n6371), .C(BIST_PATTERN[6]), .D(
        n6373), .E(AD6I), .F(n6436), .Y(n_9558) );
    zao222b U2308 ( .A(SRAM_RDATA_SEL_5), .B(n6371), .C(BIST_PATTERN[5]), .D(
        n6373), .E(AD5I), .F(n6436), .Y(n_9560) );
    zao222b U2309 ( .A(SRAM_RDATA_SEL_4), .B(n6371), .C(BIST_PATTERN[4]), .D(
        n6373), .E(AD4I), .F(n6436), .Y(n_9562) );
    zao222b U2310 ( .A(SRAM_RDATA_SEL_3), .B(n6371), .C(BIST_PATTERN[3]), .D(
        n6373), .E(AD3I), .F(n6436), .Y(n_9564) );
    zao222b U2311 ( .A(SRAM_RDATA_SEL_2), .B(n6371), .C(BIST_PATTERN[2]), .D(
        n6373), .E(AD2I), .F(n6436), .Y(n_9566) );
    zao222b U2312 ( .A(SRAM_RDATA_SEL_1), .B(n6371), .C(BIST_PATTERN[1]), .D(
        n6373), .E(AD1I), .F(n6436), .Y(n_9568) );
    zao222b U2313 ( .A(SRAM_RDATA_SEL_0), .B(n6371), .C(BIST_PATTERN[0]), .D(
        n6373), .E(AD0I), .F(n6436), .Y(n_9570) );
    zao222b U2314 ( .A(SRAM_RDATA_SEL_15), .B(n6368), .C(BIST_PATTERN[15]), 
        .D(n6369), .E(n6348), .F(AD15I), .Y(n_10216) );
    zao222b U2315 ( .A(SRAM_RDATA_SEL_14), .B(n6368), .C(BIST_PATTERN[14]), 
        .D(n6369), .E(n6348), .F(AD14I), .Y(n_10218) );
    zao222b U2316 ( .A(SRAM_RDATA_SEL_13), .B(n6368), .C(BIST_PATTERN[13]), 
        .D(n6369), .E(n6348), .F(AD13I), .Y(n_10220) );
    zao222b U2317 ( .A(SRAM_RDATA_SEL_12), .B(n6368), .C(BIST_PATTERN[12]), 
        .D(n6369), .E(n6348), .F(AD12I), .Y(n_10222) );
    zao222b U2318 ( .A(SRAM_RDATA_SEL_11), .B(n6368), .C(BIST_PATTERN[11]), 
        .D(n6369), .E(n6348), .F(AD11I), .Y(n_10224) );
    zao222b U2319 ( .A(SRAM_RDATA_SEL_10), .B(n6368), .C(BIST_PATTERN[10]), 
        .D(n6369), .E(n6348), .F(AD10I), .Y(n_10226) );
    zao222b U2320 ( .A(SRAM_RDATA_SEL_9), .B(n6368), .C(BIST_PATTERN[9]), .D(
        n6369), .E(n6348), .F(AD9I), .Y(n_10228) );
    zao222b U2321 ( .A(SRAM_RDATA_SEL_8), .B(n6368), .C(BIST_PATTERN[8]), .D(
        n6369), .E(n6348), .F(AD8I), .Y(n_10230) );
    zaoi21d U2322 ( .A(n6429), .B(n6435), .C(BIST_RUN_C), .Y(BIST_RUN4051) );
    zan2d U2323 ( .A(PM_EN), .B(n6437), .Y(DEBUG02974_2) );
    zao222b U2324 ( .A(SRAM_RDATA_SEL_23), .B(n6366), .C(BIST_PATTERN[23]), 
        .D(n6367), .E(n6342), .F(AD23I), .Y(n_10876) );
    zao222b U2325 ( .A(SRAM_RDATA_SEL_22), .B(n6366), .C(BIST_PATTERN[22]), 
        .D(n6367), .E(n6342), .F(AD22I), .Y(n_10878) );
    zao222b U2326 ( .A(SRAM_RDATA_SEL_21), .B(n6366), .C(BIST_PATTERN[21]), 
        .D(n6367), .E(n6342), .F(AD21I), .Y(n_10880) );
    zao222b U2327 ( .A(SRAM_RDATA_SEL_20), .B(n6366), .C(BIST_PATTERN[20]), 
        .D(n6367), .E(n6342), .F(AD20I), .Y(n_10882) );
    zao222b U2328 ( .A(SRAM_RDATA_SEL_19), .B(n6366), .C(BIST_PATTERN[19]), 
        .D(n6367), .E(n6342), .F(AD19I), .Y(n_10884) );
    zao222b U2329 ( .A(SRAM_RDATA_SEL_18), .B(n6366), .C(BIST_PATTERN[18]), 
        .D(n6367), .E(n6342), .F(AD18I), .Y(n_10886) );
    zao222b U2330 ( .A(SRAM_RDATA_SEL_17), .B(n6366), .C(BIST_PATTERN[17]), 
        .D(n6367), .E(n6342), .F(AD17I), .Y(n_10888) );
    zao222b U2331 ( .A(SRAM_RDATA_SEL_16), .B(n6366), .C(BIST_PATTERN[16]), 
        .D(n6367), .E(n6342), .F(AD16I), .Y(n_10890) );
    zao222b U2332 ( .A(SRAM_RDATA_SEL_31), .B(n6370), .C(BIST_PATTERN[31]), 
        .D(n6372), .E(n6353), .F(AD31I), .Y(n_11536) );
    zao222b U2333 ( .A(SRAM_RDATA_SEL_30), .B(n6370), .C(BIST_PATTERN[30]), 
        .D(n6372), .E(n6353), .F(AD30I), .Y(n_11538) );
    zao222b U2334 ( .A(SRAM_RDATA_SEL_29), .B(n6370), .C(BIST_PATTERN[29]), 
        .D(n6372), .E(n6353), .F(AD29I), .Y(n_11540) );
    zao222b U2335 ( .A(SRAM_RDATA_SEL_28), .B(n6370), .C(BIST_PATTERN[28]), 
        .D(n6372), .E(n6353), .F(AD28I), .Y(n_11542) );
    zao222b U2336 ( .A(SRAM_RDATA_SEL_27), .B(n6370), .C(BIST_PATTERN[27]), 
        .D(n6372), .E(n6353), .F(AD27I), .Y(n_11544) );
    zao222b U2337 ( .A(SRAM_RDATA_SEL_26), .B(n6370), .C(BIST_PATTERN[26]), 
        .D(n6372), .E(n6353), .F(AD26I), .Y(n_11546) );
    zao222b U2338 ( .A(SRAM_RDATA_SEL_25), .B(n6370), .C(BIST_PATTERN[25]), 
        .D(n6372), .E(n6353), .F(AD25I), .Y(n_11548) );
    zao222b U2339 ( .A(SRAM_RDATA_SEL_24), .B(n6370), .C(BIST_PATTERN[24]), 
        .D(n6372), .E(n6353), .F(AD24I), .Y(n_11550) );
    zor4b U2340 ( .A(n6438), .B(n6439), .C(n6440), .D(n6441), .Y(CFGD0) );
    zor4b U2341 ( .A(n6442), .B(n6443), .C(n6444), .D(n6445), .Y(CFGD1) );
    zor6b U2342 ( .A(n6446), .B(n6447), .C(n6448), .D(n6449), .E(n6450), .F(
        n6451), .Y(CFGD2) );
    zor4b U2343 ( .A(n6452), .B(n6453), .C(n6454), .D(n6455), .Y(CFGD3) );
    zor4b U2344 ( .A(n6456), .B(n6457), .C(n6458), .D(n6459), .Y(CFGD4) );
    zor4b U2345 ( .A(n6460), .B(n6461), .C(n6462), .D(n6463), .Y(CFGD5) );
    zor4b U2346 ( .A(n6464), .B(n6465), .C(n6466), .D(n6467), .Y(CFGD6) );
    zor3b U2347 ( .A(n6468), .B(n6469), .C(n6470), .Y(CFGD7) );
    zor5b U2348 ( .A(n6471), .B(n6472), .C(n6473), .D(n6474), .E(n6475), .Y(
        CFGD8) );
    zor4b U2349 ( .A(n6476), .B(n6477), .C(n6478), .D(n6479), .Y(CFGD9) );
    zor6b U2350 ( .A(n6480), .B(n6481), .C(n6482), .D(n6483), .E(n6484), .F(
        n6485), .Y(CFGD10) );
    zor5b U2351 ( .A(n6486), .B(n6487), .C(n6488), .D(n6489), .E(n6490), .Y(
        CFGD11) );
    zor4b U2352 ( .A(n6491), .B(n6492), .C(n6493), .D(n6494), .Y(CFGD12) );
    zor4b U2353 ( .A(n6495), .B(n6496), .C(n6497), .D(n6498), .Y(CFGD13) );
    zor4b U2354 ( .A(n6499), .B(n6500), .C(n6501), .D(n6502), .Y(CFGD14) );
    zor5b U2355 ( .A(n6503), .B(n6504), .C(n6505), .D(n6506), .E(n6507), .Y(
        CFGD15) );
    zor4b U2356 ( .A(n6508), .B(n6509), .C(n6510), .D(n6511), .Y(CFGD16) );
    zor4b U2357 ( .A(n6512), .B(n6513), .C(n6514), .D(n6515), .Y(CFGD17) );
    zor5b U2358 ( .A(n6516), .B(n6517), .C(n6518), .D(n6519), .E(n6520), .Y(
        CFGD18) );
    zor6b U2359 ( .A(n6521), .B(n6522), .C(n6523), .D(n6524), .E(n6525), .F(
        n6526), .Y(CFGD19) );
    zor5b U2360 ( .A(n6527), .B(n6528), .C(n6529), .D(n6530), .E(n6531), .Y(
        CFGD20) );
    zor5b U2361 ( .A(n6532), .B(n6533), .C(n6534), .D(n6535), .E(n6536), .Y(
        CFGD21) );
    zor5b U2362 ( .A(n6537), .B(n6538), .C(n6539), .D(n6540), .E(n6541), .Y(
        CFGD22) );
    zor4b U2363 ( .A(n6542), .B(n6543), .C(n6544), .D(n6545), .Y(CFGD23) );
    zor5b U2364 ( .A(n6546), .B(n6547), .C(n6548), .D(n6549), .E(n6550), .Y(
        CFGD24) );
    zor4b U2365 ( .A(n6551), .B(n6552), .C(n6553), .D(n6554), .Y(CFGD25) );
    zor4b U2366 ( .A(n6555), .B(n6556), .C(n6557), .D(n6558), .Y(CFGD26) );
    zor4b U2367 ( .A(n6559), .B(n6560), .C(n6561), .D(n6562), .Y(CFGD27) );
    zor6b U2368 ( .A(n6563), .B(n6564), .C(n6565), .D(n6566), .E(n6567), .F(
        n6568), .Y(CFGD28) );
    zor6b U2369 ( .A(n6569), .B(n6570), .C(n6571), .D(n6572), .E(n6573), .F(
        n6574), .Y(CFGD29) );
    zor4b U2370 ( .A(n6575), .B(n6576), .C(n6577), .D(n6578), .Y(CFGD30) );
    zor4b U2371 ( .A(n6579), .B(n6580), .C(n6581), .D(n6582), .Y(CFGD31) );
    zoa21d U2372 ( .A(AD0I), .B(AD2I), .C(AD1I), .Y(n6585) );
    zoa21d U2373 ( .A(n6587), .B(n6588), .C(TSERRS), .Y(n6412) );
    zoa21d U2374 ( .A(n6589), .B(n6588), .C(TMABORTS), .Y(n6423) );
    zoa21d U2375 ( .A(n6590), .B(n6588), .C(TTABORTR), .Y(n6413) );
    zor3b U2376 ( .A(n6609), .B(n6608), .C(n6607), .Y(n6610) );
    zor2d U2377 ( .A(n6613), .B(n7134), .Y(n6617) );
    zivh U2378 ( .A(AD2I), .Y(n6620) );
    zivh U2379 ( .A(AD3I), .Y(n6622) );
    zivh U2380 ( .A(AD4I), .Y(n6624) );
    zivh U2381 ( .A(AD7I), .Y(n6630) );
    zor2d U2382 ( .A(CBE1I_), .B(n6612), .Y(n6632) );
    zor3b U2383 ( .A(n6608), .B(n6609), .C(n6644), .Y(n6645) );
    zor2d U2384 ( .A(CBE3I_), .B(n6612), .Y(n6646) );
    zor2d U2385 ( .A(CBE2I_), .B(n6612), .Y(n6661) );
    zor3b U2386 ( .A(PA4I), .B(n6608), .C(n6644), .Y(n6700) );
    zor2d U2387 ( .A(n6613), .B(n6729), .Y(n6730) );
    zor4b U2388 ( .A(SLAVEMODE), .B(BIST_RUN), .C(SLAVE_ACT), .D(n6743), .Y(
        n6764) );
    zor3b U2389 ( .A(PA4I), .B(PA6I), .C(n6607), .Y(n6766) );
    zor4b U2390 ( .A(n6609), .B(n6813), .C(n6606), .D(n6608), .Y(n6814) );
    zor4b U2391 ( .A(PA5I), .B(n6813), .C(PA4I), .D(PA6I), .Y(n6824) );
    zor3b U2392 ( .A(PA4I), .B(n6608), .C(n6607), .Y(n6825) );
    zor3b U2393 ( .A(PA4I), .B(PA6I), .C(n6644), .Y(n6878) );
    zor3b U2394 ( .A(PA6I), .B(n6609), .C(n6644), .Y(n6880) );
    zor3b U2395 ( .A(PA6I), .B(n6609), .C(n6607), .Y(n6922) );
    zor3b U2396 ( .A(FUNCSEL[1]), .B(FUNCSEL[0]), .C(n7021), .Y(n7022) );
    zmux21ld U2397 ( .A(n6636), .B(n6618), .S(n7045), .Y(n_8054) );
    zmux21ld U2398 ( .A(n6638), .B(n6619), .S(n7045), .Y(n_8052) );
    zmux21ld U2399 ( .A(n6639), .B(n6620), .S(n7045), .Y(n_8050) );
    zmux21ld U2400 ( .A(n6640), .B(n6622), .S(n7045), .Y(n_8048) );
    zmux21ld U2401 ( .A(n6641), .B(n6624), .S(n7045), .Y(n_8046) );
    zmux21ld U2402 ( .A(n6642), .B(n6626), .S(n7045), .Y(n_8044) );
    zmux21ld U2403 ( .A(n6643), .B(n6628), .S(n7045), .Y(n_8042) );
    zmux21ld U2404 ( .A(n6604), .B(n6630), .S(n7045), .Y(n_8040) );
    zmux21ld U2405 ( .A(n6693), .B(n6620), .S(n7046), .Y(n_5142) );
    zmux21ld U2406 ( .A(n6694), .B(n6622), .S(n7046), .Y(n_5140) );
    zmux21ld U2407 ( .A(n6695), .B(n6624), .S(n7046), .Y(n_5138) );
    zmux21ld U2408 ( .A(n6696), .B(n6626), .S(n7046), .Y(n_5136) );
    zmux21ld U2409 ( .A(n6697), .B(n6628), .S(n7046), .Y(n_5134) );
    zmux21ld U2410 ( .A(n6698), .B(n6630), .S(n7046), .Y(n_5132) );
    zmux21ld U2411 ( .A(n6731), .B(n6622), .S(n7047), .Y(TrkSpd3743_1) );
    zmux21ld U2412 ( .A(n6732), .B(n6620), .S(n7047), .Y(TrkSpd3743_0) );
    zmux21ld U2413 ( .A(n6776), .B(n6630), .S(n6376), .Y(SUBVID02822_7) );
    zmux21ld U2414 ( .A(n6777), .B(n6628), .S(n6376), .Y(SUBVID02822_6) );
    zmux21ld U2415 ( .A(n6778), .B(n6626), .S(n6376), .Y(SUBVID02822_5) );
    zmux21ld U2416 ( .A(n6779), .B(n6624), .S(n6376), .Y(SUBVID02822_4) );
    zmux21ld U2417 ( .A(n6780), .B(n6622), .S(n6376), .Y(SUBVID02822_3) );
    zmux21ld U2418 ( .A(n6781), .B(n6620), .S(n6376), .Y(SUBVID02822_2) );
    zmux21ld U2419 ( .A(n6782), .B(n6619), .S(n6376), .Y(SUBVID02822_1) );
    zmux21ld U2420 ( .A(n6783), .B(n6618), .S(n6376), .Y(SUBVID02822_0) );
    zmux21ld U2421 ( .A(n6810), .B(n6628), .S(n7047), .Y(RxDataDly3781_2) );
    zmux21ld U2422 ( .A(n6811), .B(n6626), .S(n7047), .Y(RxDataDly3781_1) );
    zmux21ld U2423 ( .A(n6812), .B(n6624), .S(n7047), .Y(RxDataDly3781_0) );
    zmux21ld U2424 ( .A(n6869), .B(n6630), .S(n7049), .Y(PHYOPT13477_7) );
    zmux21ld U2425 ( .A(n6870), .B(n6628), .S(n7049), .Y(PHYOPT13477_6) );
    zmux21ld U2426 ( .A(n6871), .B(n6626), .S(n7049), .Y(PHYOPT13477_5) );
    zmux21ld U2427 ( .A(n6872), .B(n6624), .S(n7049), .Y(PHYOPT13477_4) );
    zmux21ld U2428 ( .A(n6873), .B(n6622), .S(n7049), .Y(PHYOPT13477_3) );
    zmux21ld U2429 ( .A(n6874), .B(n6620), .S(n7049), .Y(PHYOPT13477_2) );
    zmux21ld U2430 ( .A(n6875), .B(n6619), .S(n7049), .Y(PHYOPT13477_1) );
    zmux21ld U2431 ( .A(n6876), .B(n6618), .S(n7049), .Y(PHYOPT13477_0) );
    zmux21ld U2432 ( .A(n6746), .B(n6630), .S(n7050), .Y(PHYMON_EN_H4404) );
    zmux21ld U2433 ( .A(n6747), .B(n6628), .S(n7050), .Y(PHYMON_EN_G4398) );
    zmux21ld U2434 ( .A(n6748), .B(n6626), .S(n7050), .Y(PHYMON_EN_F4392) );
    zmux21ld U2435 ( .A(n6749), .B(n6624), .S(n7050), .Y(PHYMON_EN_E4386) );
    zmux21ld U2436 ( .A(n6750), .B(n6622), .S(n7050), .Y(PHYMON_EN_D4380) );
    zmux21ld U2437 ( .A(n6752), .B(n6620), .S(n7050), .Y(PHYMON_EN_C4374) );
    zmux21ld U2438 ( .A(n6754), .B(n6619), .S(n7050), .Y(PHYMON_EN_B4368) );
    zmux21ld U2439 ( .A(n6756), .B(n6618), .S(n7050), .Y(PHYMON_EN_A4362) );
    zmux21ld U2440 ( .A(n6884), .B(n6624), .S(n6381), .Y(MWRMEN2052) );
    zmux21ld U2441 ( .A(n6885), .B(n6619), .S(n6381), .Y(MMSPACE2040) );
    zmux21ld U2442 ( .A(n6886), .B(n6619), .S(n7047), .Y(LockSpd3705_1) );
    zmux21ld U2443 ( .A(n6887), .B(n6618), .S(n7047), .Y(LockSpd3705_0) );
    zmux21ld U2444 ( .A(n6896), .B(n6618), .S(n6381), .Y(IOSPACE2034) );
    zmux21ld U2445 ( .A(n6723), .B(n6630), .S(n7051), .Y(INTLN2337_7) );
    zmux21ld U2446 ( .A(n6722), .B(n6628), .S(n7051), .Y(INTLN2337_6) );
    zmux21ld U2447 ( .A(n6724), .B(n6626), .S(n7051), .Y(INTLN2337_5) );
    zmux21ld U2448 ( .A(n6721), .B(n6624), .S(n7051), .Y(INTLN2337_4) );
    zmux21ld U2449 ( .A(n6725), .B(n6622), .S(n7051), .Y(INTLN2337_3) );
    zmux21ld U2450 ( .A(n6726), .B(n6620), .S(n7051), .Y(INTLN2337_2) );
    zmux21ld U2451 ( .A(n6727), .B(n6619), .S(n7051), .Y(INTLN2337_1) );
    zmux21ld U2452 ( .A(n6728), .B(n6618), .S(n7051), .Y(INTLN2337_0) );
    zmux21ld U2453 ( .A(n6923), .B(n6630), .S(n7047), .Y(FastStart3819) );
    zmux21ld U2454 ( .A(n6959), .B(n6630), .S(n7052), .Y(DEBUGC3325_7) );
    zmux21ld U2455 ( .A(n6960), .B(n6628), .S(n7052), .Y(DEBUGC3325_6) );
    zmux21ld U2456 ( .A(n6961), .B(n6626), .S(n7052), .Y(DEBUGC3325_5) );
    zmux21ld U2457 ( .A(n6962), .B(n6624), .S(n7052), .Y(DEBUGC3325_4) );
    zmux21ld U2458 ( .A(n6963), .B(n6622), .S(n7052), .Y(DEBUGC3325_3) );
    zmux21ld U2459 ( .A(n6964), .B(n6620), .S(n7052), .Y(DEBUGC3325_2) );
    zmux21ld U2460 ( .A(n6965), .B(n6619), .S(n7052), .Y(DEBUGC3325_1) );
    zmux21ld U2461 ( .A(n6966), .B(n6618), .S(n7052), .Y(DEBUGC3325_0) );
    zmux21ld U2462 ( .A(n6983), .B(n6630), .S(n7054), .Y(DEBUG83126_7) );
    zmux21ld U2463 ( .A(n6984), .B(n6628), .S(n7054), .Y(DEBUG83126_6) );
    zmux21ld U2464 ( .A(n6985), .B(n6626), .S(n7054), .Y(DEBUG83126_5) );
    zmux21ld U2465 ( .A(n6986), .B(n6624), .S(n7054), .Y(DEBUG83126_4) );
    zmux21ld U2466 ( .A(n6987), .B(n6622), .S(n7054), .Y(DEBUG83126_3) );
    zmux21ld U2467 ( .A(n6988), .B(n6620), .S(n7054), .Y(DEBUG83126_2) );
    zmux21ld U2468 ( .A(n6989), .B(n6619), .S(n7054), .Y(DEBUG83126_1) );
    zmux21ld U2469 ( .A(n6990), .B(n6618), .S(n7054), .Y(DEBUG83126_0) );
    zmux21ld U2470 ( .A(n7013), .B(n6630), .S(n7055), .Y(DEBUG02974_7) );
    zmux21ld U2471 ( .A(n7014), .B(n6628), .S(n7055), .Y(DEBUG02974_6) );
    zmux21ld U2472 ( .A(n7015), .B(n6626), .S(n7055), .Y(DEBUG02974_5) );
    zmux21ld U2473 ( .A(n7016), .B(n6624), .S(n7055), .Y(DEBUG02974_4) );
    zmux21ld U2474 ( .A(n7017), .B(n6622), .S(n7055), .Y(DEBUG02974_3) );
    zmux21ld U2475 ( .A(FCFG), .B(n6619), .S(n7055), .Y(DEBUG02974_1) );
    zmux21ld U2476 ( .A(n7019), .B(n6618), .S(n7055), .Y(DEBUG02974_0) );
    zmux21ld U2477 ( .A(n7027), .B(n6630), .S(n7056), .Y(CACHLN72206) );
    zmux21ld U2478 ( .A(n7028), .B(n6628), .S(n7056), .Y(CACHLN62200) );
    zmux21ld U2479 ( .A(n7029), .B(n6626), .S(n7056), .Y(CACHLN52194) );
    zmux21ld U2480 ( .A(n7030), .B(n6624), .S(n7056), .Y(CACHLN42188) );
    zmux21ld U2481 ( .A(n7033), .B(n6622), .S(n7056), .Y(CACHLN32182) );
    zmux21ld U2482 ( .A(n7040), .B(n6620), .S(n7056), .Y(CACHLN22176) );
    zmux21ld U2483 ( .A(n7042), .B(n6619), .S(n7056), .Y(CACHLN12170) );
    zmux21ld U2484 ( .A(n7043), .B(n6618), .S(n7056), .Y(CACHLN02164) );
    zmux21ld U2485 ( .A(n7041), .B(n6620), .S(n6381), .Y(BMASTREN2046) );
    zmux21ld U2486 ( .A(n7025), .B(n6618), .S(n6418), .Y(BACK_EN5715) );
    zao222b U2487 ( .A(IOBA9), .B(n6586), .C(FLADJ1), .D(n6416), .E(USBLEGSUP
        [9]), .F(n6390), .Y(n7057) );
    zao211b U2488 ( .A(USBLEGCTLSTS[9]), .B(n7125), .C(n6364), .D(n7057), .Y(
        n6478) );
    zao211b U2489 ( .A(PME_EN), .B(n6362), .C(n6360), .D(n6364), .Y(n6473) );
    zao222b U2490 ( .A(REVID_BACK_0), .B(n7058), .C(BIST_PATTERN[8]), .D(n7059
        ), .E(UIRQACT), .F(n7060), .Y(n6471) );
    zao222b U2491 ( .A(n6391), .B(TMOUT_PARM[0]), .C(n6361), .D(SUBVID1_0), 
        .E(DEBUG9_0), .F(n7063), .Y(n7061) );
    zao222b U2492 ( .A(n7068), .B(LAT_TM_0), .C(CTRL_F[0]), .D(n7069), .E(
        BypassDiv4), .F(n7070), .Y(n7067) );
    zor4b U2493 ( .A(n7067), .B(n7071), .C(n7061), .D(n7064), .Y(n6475) );
    zao222b U2494 ( .A(n7074), .B(n7075), .C(n7037), .D(n7076), .E(
        USBLEGCTLSTS[7]), .F(n6389), .Y(n7073) );
    zao211b U2495 ( .A(USBLEGSUP[7]), .B(n6422), .C(n7073), .D(n7077), .Y(
        n6470) );
    zao211b U2496 ( .A(n6374), .B(REVID_BACK_5), .C(n7078), .D(n7079), .Y(
        n6462) );
    zao222b U2497 ( .A(USBLEGCTLSTS[4]), .B(n6389), .C(n7037), .D(n7080), .E(
        USBLEGSUP[4]), .F(n6390), .Y(n6456) );
    zao222b U2498 ( .A(SRAM_ADDR[4]), .B(n7072), .C(MWRMEN), .D(n7083), .E(
        n6393), .F(INTLN_4), .Y(n7082) );
    zao211b U2499 ( .A(n7066), .B(PHYMON_EN_E), .C(n7082), .D(n7081), .Y(n6459
        ) );
    zao211b U2500 ( .A(USBLEGCTLSTS[31]), .B(n7125), .C(n6365), .D(n7085), .Y(
        n6581) );
    zao222b U2501 ( .A(DEBUGF_7), .B(n6593), .C(DIS_TERM_ON_H), .D(n7060), .E(
        CTRL_A[3]), .F(n7070), .Y(n6580) );
    zao211b U2502 ( .A(USBLEGCTLSTS[30]), .B(n7125), .C(n7036), .D(n7086), .Y(
        n6577) );
    zao211b U2503 ( .A(n6374), .B(REVID_BACK_3), .C(n7087), .D(n7088), .Y(
        n6454) );
    zor3b U2504 ( .A(n6363), .B(n7036), .C(n6360), .Y(n7089) );
    zao211b U2505 ( .A(USBLEGSUP[29]), .B(n6422), .C(n6591), .D(n7089), .Y(
        n6574) );
    zao222b U2506 ( .A(MAXLAT5), .B(n7084), .C(BIST_PATTERN[29]), .D(n7059), 
        .E(SL_ERROFFSET[5]), .F(n7062), .Y(n6572) );
    zao222b U2507 ( .A(SUBSID1_5), .B(n6361), .C(Disconnect_H), .D(n6387), .E(
        SLEEPTIME_SEL), .F(n7063), .Y(n6569) );
    zao211b U2508 ( .A(USBLEGCTLSTS[28]), .B(n7125), .C(n6360), .D(n7036), .Y(
        n6566) );
    zao222b U2509 ( .A(SUBSID1_4), .B(n6361), .C(n7069), .D(TERMON_H), .E(
        DIS_SOF_RUN), .F(n7063), .Y(n6563) );
    zao211b U2510 ( .A(DIS_TERM_ON_D), .B(n7060), .C(n6592), .D(n7035), .Y(
        n6560) );
    zao211b U2511 ( .A(DIS_TERM_ON_C), .B(n7060), .C(n6594), .D(n7035), .Y(
        n6556) );
    zao211b U2512 ( .A(USBLEGCTLSTS[25]), .B(n7125), .C(n7090), .D(n7091), .Y(
        n6553) );
    zor4b U2513 ( .A(n6360), .B(n6365), .C(n6595), .D(n7092), .Y(n6549) );
    zao222b U2514 ( .A(IOBA24), .B(n6586), .C(n7066), .D(TERMON_E), .E(
        TURN_PARM[0]), .F(n7063), .Y(n6546) );
    zao222b U2515 ( .A(REVID7), .B(n7058), .C(n7068), .D(n7095), .E(n7093), 
        .F(n6416), .Y(n7094) );
    zao222b U2516 ( .A(SUBSID0_7), .B(n6361), .C(MINGNT7), .D(n7084), .E(
        SLAVE_ERR), .F(n7062), .Y(n7097) );
    zor5b U2517 ( .A(n6363), .B(n6365), .C(n7094), .D(n7097), .E(n7096), .Y(
        n6545) );
    zao211b U2518 ( .A(REVID6), .B(n7058), .C(n6365), .D(n6596), .Y(n6537) );
    zao211b U2519 ( .A(REVID5), .B(n7058), .C(n6363), .D(n6597), .Y(n6532) );
    zao211b U2520 ( .A(REVID4), .B(n7058), .C(n7083), .D(n6598), .Y(n6527) );
    zao211b U2521 ( .A(n6374), .B(REVID_BACK_2), .C(n6360), .D(n6599), .Y(
        n6449) );
    zao222b U2522 ( .A(BIST_PATTERN[2]), .B(n7059), .C(sync_jend), .D(n6593), 
        .E(SOF_DISCONN_CHK), .F(n7070), .Y(n6448) );
    zao222b U2523 ( .A(REVID3), .B(n7058), .C(n7098), .D(n6416), .E(
        USBLEGCTLSTS[19]), .F(n6425), .Y(n6524) );
    zao222b U2524 ( .A(IOBA19), .B(n6586), .C(BIST_PATTERN[19]), .D(n7059), 
        .E(n7066), .F(RxData_C), .Y(n6521) );
    zao211b U2525 ( .A(REVID2), .B(n7058), .C(n6360), .D(n6600), .Y(n6516) );
    zao211b U2526 ( .A(USBLEGCTLSTS[17]), .B(n7125), .C(n7099), .D(n7100), .Y(
        n6514) );
    zao211b U2527 ( .A(CTRL_D[1]), .B(n7070), .C(n7035), .D(n7101), .Y(n6513)
         );
    zao211b U2528 ( .A(USBLEGCTLSTS[16]), .B(n7125), .C(n7102), .D(n7103), .Y(
        n6510) );
    zao222b U2529 ( .A(BIST_PATTERN[15]), .B(n7059), .C(IOBA15), .D(n6586), 
        .E(USBLEGSUP[15]), .F(n7124), .Y(n6503) );
    zao222b U2530 ( .A(DEBUGD_6), .B(n6593), .C(n7068), .D(LAT_TM_6), .E(
        DISPRST), .F(n7060), .Y(n6500) );
    zao222b U2531 ( .A(IOBA13), .B(n6586), .C(FLADJ5), .D(n6416), .E(USBLEGSUP
        [13]), .F(n6390), .Y(n7104) );
    zao211b U2532 ( .A(USBLEGCTLSTS[13]), .B(n7125), .C(n7037), .D(n7104), .Y(
        n6497) );
    zao222b U2533 ( .A(IOBA12), .B(n6586), .C(FLADJ4), .D(n6416), .E(USBLEGSUP
        [12]), .F(n7124), .Y(n7105) );
    zao211b U2534 ( .A(USBLEGCTLSTS[12]), .B(n7125), .C(n6360), .D(n7105), .Y(
        n6493) );
    zao222b U2535 ( .A(BIST_PATTERN[11]), .B(n7059), .C(IOBA11), .D(n6586), 
        .E(USBLEGSUP[11]), .F(n7124), .Y(n6486) );
    zao222b U2536 ( .A(IOBA10), .B(n6586), .C(FLADJ2), .D(n6416), .E(USBLEGSUP
        [10]), .F(n6390), .Y(n6483) );
    zao222b U2537 ( .A(n7066), .B(Squelch_A), .C(n6361), .D(SUBVID1_2), .E(
        SLQUEUEADDR[10]), .F(n7065), .Y(n6480) );
    zao211b U2538 ( .A(n6374), .B(REVID_BACK_1), .C(n6360), .D(n6363), .Y(
        n7106) );
    zao222b U2539 ( .A(CACHLN1), .B(n7068), .C(n6361), .D(SUBVID0_1), .E(
        USBLEGSUP[1]), .F(n7124), .Y(n7108) );
    zor4b U2540 ( .A(n7108), .B(n7109), .C(n7106), .D(n7107), .Y(n6445) );
    zao222b U2541 ( .A(SRAM_ADDR[1]), .B(n7072), .C(LockSpd[1]), .D(n7069), 
        .E(EN_CHKTOGCRC), .F(n7063), .Y(n6442) );
    zao211b U2542 ( .A(n6374), .B(REVID_BACK_0), .C(n7036), .D(n6601), .Y(
        n7110) );
    zao222b U2543 ( .A(CACHLN0), .B(n7068), .C(USBLEGSUP[0]), .D(n6422), .E(
        DEBUG0_0), .F(n7060), .Y(n7112) );
    zor4b U2544 ( .A(n7112), .B(n7113), .C(n7110), .D(n7111), .Y(n6441) );
    zao222b U2545 ( .A(LockSpd[0]), .B(n7069), .C(IOSPACE), .D(n7083), .E(
        HsEnFB_Dis), .F(n7063), .Y(n6438) );
    zoa22d U2546 ( .A(n6622), .B(n6742), .C(BIST_ERR_S), .D(BIST_ERROR), .Y(
        n6434) );
    zor2d U2547 ( .A(n6613), .B(n6635), .Y(n7114) );
    zivh U2548 ( .A(n7114), .Y(n7045) );
    zor2d U2549 ( .A(n6613), .B(n6844), .Y(n7116) );
    zivh U2550 ( .A(n7116), .Y(n7049) );
    zor2d U2551 ( .A(n6613), .B(n7128), .Y(n6437) );
    zor4b U2552 ( .A(AD0I), .B(AD1I), .C(n6620), .D(n6764), .Y(n6435) );
    zor2d U2553 ( .A(n6730), .B(n6878), .Y(n7117) );
    zivh U2554 ( .A(n7117), .Y(n7056) );
    zor2d U2555 ( .A(n6730), .B(n6922), .Y(n7118) );
    zivh U2556 ( .A(n7118), .Y(n7051) );
    zor2d U2557 ( .A(n6613), .B(n7132), .Y(n7119) );
    zivh U2558 ( .A(n7119), .Y(n7054) );
    zor2d U2559 ( .A(n6645), .B(n6730), .Y(n7120) );
    zivh U2560 ( .A(n7120), .Y(n7047) );
    zor2d U2561 ( .A(n6613), .B(n6647), .Y(n7121) );
    zivh U2562 ( .A(n7121), .Y(n7046) );
    zor2d U2563 ( .A(n6700), .B(n6730), .Y(n7122) );
    zivh U2564 ( .A(n7122), .Y(n7052) );
    zor2d U2565 ( .A(n6613), .B(n7126), .Y(n7123) );
    zivh U2566 ( .A(n7123), .Y(n7050) );
    zivh U2567 ( .A(n6632), .Y(n6426) );
    zivh U2568 ( .A(n6661), .Y(n6417) );
    zor4b U2569 ( .A(n6723), .B(n6724), .C(n6721), .D(n6722), .Y(n6421) );
    zor3b U2570 ( .A(n7021), .B(n7038), .C(n7039), .Y(n7095) );
endmodule


module HS_DBG_OPREG ( ADI, EN_DBG_PORT, DBGPORT_R00G, DBGPORT_R01G, 
    DBGPORT_R02G, DBGPORT_R03G, DBGPORT_R04G, DBGPORT_R05G, DBGPORT_R10G, 
    DBGPORT_R11G, DBGPORT_SC, DBGPORT_PID, DBGPORT_ADDR, DBG_COMPL, 
    DBG_XACTERR, PORT_ENDIS, PORT_SUSPEND, PORT_RESET, DBG_RXBCNT, DBG_RXPID, 
    DBG_ENABLE_WC, PCICLK, PCICLK_FREE, CMDRST_ );
input  [31:0] ADI;
input  [3:0] DBG_RXBCNT;
output [31:0] DBGPORT_SC;
input  [7:0] DBG_RXPID;
output [31:0] DBGPORT_PID;
output [31:0] DBGPORT_ADDR;
input  EN_DBG_PORT, DBGPORT_R00G, DBGPORT_R01G, DBGPORT_R02G, DBGPORT_R03G, 
    DBGPORT_R04G, DBGPORT_R05G, DBGPORT_R10G, DBGPORT_R11G, DBG_COMPL, 
    DBG_XACTERR, PORT_ENDIS, PORT_SUSPEND, PORT_RESET, PCICLK, PCICLK_FREE, 
    CMDRST_;
output DBG_ENABLE_WC;
    wire DBG_DONE, DBG_LENGTH484_3, SPAREO6, DBG_RCVPID572_1, DBG_TXPID_3, 
        DBG_ERRGD, DBG_LENGTH_3, DBG_TOKEN648_0, DBG_TOKEN_0, DBG_TXPID610_7, 
        DBG_RCVPID_4, PORT_BLOCK, DBG_ADDR722_0, DBG_WR, DBG_ADDR_0, DBG_WR403, 
        DBG_ENDP_1, DBG_RCVPID_3, SPAREO0_, DBG_ENDP760_2, DBG_TXPID610_0, 
        DBG_TOKEN_7, DBG_TOKEN648_7, DBG_TXPID_4, DBG_RCVPID572_6, SPAREO1, 
        DBG_TXPID610_1, SPAREO9, DBG_ENDP760_3, DBG_ENDP_0, DBG_RCVPID_2, 
        DBG_ADDR722_6, DBG_ADDR_6, SPAREO0, DBG_TXPID_5, DBG_RCVPID572_7, 
        DBG_TOKEN648_6, DBG_TOKEN_6, DBG_TOKEN648_1, DBG_OWNER141, DBG_TOKEN_1, 
        DBG_TXPID_2, DBG_RCVPID572_0, DBG_LENGTH_2, SPAREO7, DBG_LENGTH484_2, 
        DBG_ADDR722_1, DBG_ERRGD289, DBG_ADDR_1, DBG_RCVPID_5, DBG_TXPID610_6, 
        DBG_LENGTH484_0, DBG_ENABLE178, SPAREO5, DBG_OWNER, DBG_LENGTH_0, 
        DBG_TXPID_0, DBG_GO, DBG_RCVPID572_2, DBG_TOKEN_3, DBG_TOKEN648_3, 
        DBG_DONE215, DBG_TXPID610_4, DBG_GO366, DBG_RCVPID_7, PORT_BLOCK_T326, 
        DBG_ADDR_3, DBG_ADDR722_3, DBG_ADDR_4, DBG_ADDR722_4, DBG_RCVPID_0, 
        DBG_ENDP_2, DBG_ENDP760_1, DBG_TXPID610_3, PORT_BLOCK_T, DBG_TOKEN_4, 
        DBG_TOKEN648_4, DBG_RCVPID572_5, DBG_TXPID_7, SPAREO2, DBG_TXPID610_2, 
        DBG_ENDP760_0, DBG_RCVPID_1, DBG_ENDP_3, DBG_ADDR_5, DBG_ADDR722_5, 
        SPAREO3, SPAREO1_, DBG_RCVPID572_4, DBG_TXPID_6, DBG_TOKEN_5, 
        DBG_TOKEN648_5, DBG_TOKEN_2, DBG_LENGTH_1, DBG_TOKEN648_2, DBG_TXPID_1, 
        DBG_RCVPID572_3, SPAREO4, DBG_LENGTH484_1, DBG_INUSE252, DBG_INUSE, 
        DBG_ADDR_2, DBG_ADDR722_2, DBG_RCVPID_6, a425, DBG_ENABLE, 
        DBG_TXPID610_5, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
        n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
        n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
        n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
        n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
        n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, 
        n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089;
    assign DBGPORT_SC[31] = 1'b0;
    assign DBGPORT_SC[29] = 1'b0;
    assign DBGPORT_SC[27] = 1'b0;
    assign DBGPORT_SC[26] = 1'b0;
    assign DBGPORT_SC[25] = 1'b0;
    assign DBGPORT_SC[24] = 1'b0;
    assign DBGPORT_SC[23] = 1'b0;
    assign DBGPORT_SC[22] = 1'b0;
    assign DBGPORT_SC[21] = 1'b0;
    assign DBGPORT_SC[20] = 1'b0;
    assign DBGPORT_SC[19] = 1'b0;
    assign DBGPORT_SC[18] = 1'b0;
    assign DBGPORT_SC[17] = 1'b0;
    assign DBGPORT_SC[15] = 1'b0;
    assign DBGPORT_SC[14] = 1'b0;
    assign DBGPORT_SC[13] = 1'b0;
    assign DBGPORT_SC[12] = 1'b0;
    assign DBGPORT_SC[11] = 1'b0;
    assign DBGPORT_SC[9] = 1'b0;
    assign DBGPORT_PID[31] = 1'b0;
    assign DBGPORT_PID[30] = 1'b0;
    assign DBGPORT_PID[29] = 1'b0;
    assign DBGPORT_PID[28] = 1'b0;
    assign DBGPORT_PID[27] = 1'b0;
    assign DBGPORT_PID[26] = 1'b0;
    assign DBGPORT_PID[25] = 1'b0;
    assign DBGPORT_PID[24] = 1'b0;
    assign DBGPORT_ADDR[31] = 1'b0;
    assign DBGPORT_ADDR[30] = 1'b0;
    assign DBGPORT_ADDR[29] = 1'b0;
    assign DBGPORT_ADDR[28] = 1'b0;
    assign DBGPORT_ADDR[27] = 1'b0;
    assign DBGPORT_ADDR[26] = 1'b0;
    assign DBGPORT_ADDR[25] = 1'b0;
    assign DBGPORT_ADDR[24] = 1'b0;
    assign DBGPORT_ADDR[23] = 1'b0;
    assign DBGPORT_ADDR[22] = 1'b0;
    assign DBGPORT_ADDR[21] = 1'b0;
    assign DBGPORT_ADDR[20] = 1'b0;
    assign DBGPORT_ADDR[19] = 1'b0;
    assign DBGPORT_ADDR[18] = 1'b0;
    assign DBGPORT_ADDR[17] = 1'b0;
    assign DBGPORT_ADDR[16] = 1'b0;
    assign DBGPORT_ADDR[15] = 1'b0;
    assign DBGPORT_ADDR[7] = 1'b0;
    assign DBGPORT_ADDR[6] = 1'b0;
    assign DBGPORT_ADDR[5] = 1'b0;
    assign DBGPORT_ADDR[4] = 1'b0;
    znd3b SPARE_DBG9 ( .A(SPAREO3), .B(SPAREO6), .C(1'b0), .Y(SPAREO7) );
    zdffrb SPARE_DBG0 ( .CK(PCICLK), .D(1'b0), .R(n1089), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE_DBG7 ( .A(SPAREO4), .Y(SPAREO5) );
    znr3b SPARE_DBG6 ( .A(SPAREO2), .B(PORT_BLOCK), .C(SPAREO0_), .Y(SPAREO4)
         );
    zivb SPARE_DBG8 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE_DBG1 ( .CK(PCICLK), .D(SPAREO7), .R(n1089), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zaoi211b SPARE_DBG3 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0) );
    zoai21b SPARE_DBG4 ( .A(SPAREO0), .B(n1026), .C(1'b0), .Y(SPAREO9) );
    zoai21b SPARE_DBG5 ( .A(SPAREO1), .B(n1025), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE_DBG2 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    znr2b U338 ( .A(ADI[1]), .B(ADI[0]), .Y(n1029) );
    zor2b U339 ( .A(ADI[3]), .B(a425), .Y(n1037) );
    zan2b U340 ( .A(DBGPORT_R00G), .B(ADI[2]), .Y(n1035) );
    zivb U341 ( .A(a425), .Y(n1036) );
    zaoi21b U342 ( .A(n1029), .B(n1054), .C(n1083), .Y(a425) );
    zmux21hb U343 ( .A(DBG_RCVPID_7), .B(DBG_RXPID[7]), .S(DBG_COMPL), .Y(
        DBG_RCVPID572_7) );
    zmux21hb U344 ( .A(DBG_RCVPID_6), .B(DBG_RXPID[6]), .S(DBG_COMPL), .Y(
        DBG_RCVPID572_6) );
    zmux21hb U345 ( .A(DBG_RCVPID_5), .B(DBG_RXPID[5]), .S(DBG_COMPL), .Y(
        DBG_RCVPID572_5) );
    zmux21hb U346 ( .A(DBG_RCVPID_4), .B(DBG_RXPID[4]), .S(DBG_COMPL), .Y(
        DBG_RCVPID572_4) );
    zmux21hb U347 ( .A(DBG_RCVPID_3), .B(DBG_RXPID[3]), .S(DBG_COMPL), .Y(
        DBG_RCVPID572_3) );
    zmux21hb U348 ( .A(DBG_RCVPID_2), .B(DBG_RXPID[2]), .S(DBG_COMPL), .Y(
        DBG_RCVPID572_2) );
    zmux21hb U349 ( .A(DBG_RCVPID_1), .B(DBG_RXPID[1]), .S(DBG_COMPL), .Y(
        DBG_RCVPID572_1) );
    zmux21hb U350 ( .A(DBG_RCVPID_0), .B(DBG_RXPID[0]), .S(DBG_COMPL), .Y(
        DBG_RCVPID572_0) );
    zmux21hb U351 ( .A(DBG_TXPID_7), .B(ADI[15]), .S(DBGPORT_R05G), .Y(
        DBG_TXPID610_7) );
    zmux21lb U352 ( .A(n1043), .B(n1076), .S(DBGPORT_R05G), .Y(DBG_TXPID610_6)
         );
    zmux21lb U353 ( .A(n1044), .B(n1077), .S(DBGPORT_R05G), .Y(DBG_TXPID610_5)
         );
    zmux21lb U354 ( .A(n1045), .B(n1078), .S(DBGPORT_R05G), .Y(DBG_TXPID610_4)
         );
    zmux21lb U355 ( .A(n1046), .B(n1079), .S(DBGPORT_R05G), .Y(DBG_TXPID610_3)
         );
    zmux21lb U356 ( .A(n1047), .B(n1080), .S(DBGPORT_R05G), .Y(DBG_TXPID610_2)
         );
    zmux21lb U357 ( .A(n1048), .B(n1081), .S(DBGPORT_R05G), .Y(DBG_TXPID610_1)
         );
    zmux21lb U358 ( .A(n1049), .B(n1082), .S(DBGPORT_R05G), .Y(DBG_TXPID610_0)
         );
    zmux21hb U359 ( .A(DBG_TOKEN_7), .B(ADI[7]), .S(DBGPORT_R04G), .Y(
        DBG_TOKEN648_7) );
    zmux21hb U360 ( .A(DBG_TOKEN_6), .B(ADI[6]), .S(DBGPORT_R04G), .Y(
        DBG_TOKEN648_6) );
    zmux21lb U361 ( .A(n1051), .B(n1050), .S(DBGPORT_R04G), .Y(DBG_TOKEN648_5)
         );
    zmux21lb U362 ( .A(n1052), .B(n1075), .S(DBGPORT_R04G), .Y(DBG_TOKEN648_4)
         );
    zmux21lb U363 ( .A(n1053), .B(n1083), .S(DBGPORT_R04G), .Y(DBG_TOKEN648_3)
         );
    zmux21lb U364 ( .A(n1055), .B(n1054), .S(DBGPORT_R04G), .Y(DBG_TOKEN648_2)
         );
    zmux21lb U365 ( .A(n1056), .B(n1040), .S(DBGPORT_R04G), .Y(DBG_TOKEN648_1)
         );
    zmux21lb U366 ( .A(n1057), .B(n1041), .S(DBGPORT_R04G), .Y(DBG_TOKEN648_0)
         );
    zmux21lb U367 ( .A(n1066), .B(n1076), .S(DBGPORT_R11G), .Y(DBG_ADDR722_6)
         );
    zivb U368 ( .A(ADI[14]), .Y(n1076) );
    zmux21lb U369 ( .A(n1067), .B(n1077), .S(DBGPORT_R11G), .Y(DBG_ADDR722_5)
         );
    zivb U370 ( .A(ADI[13]), .Y(n1077) );
    zmux21lb U371 ( .A(n1068), .B(n1078), .S(DBGPORT_R11G), .Y(DBG_ADDR722_4)
         );
    zivb U372 ( .A(ADI[12]), .Y(n1078) );
    zmux21lb U373 ( .A(n1069), .B(n1079), .S(DBGPORT_R11G), .Y(DBG_ADDR722_3)
         );
    zivb U374 ( .A(ADI[11]), .Y(n1079) );
    zmux21lb U375 ( .A(n1070), .B(n1080), .S(DBGPORT_R11G), .Y(DBG_ADDR722_2)
         );
    zmux21lb U376 ( .A(n1071), .B(n1081), .S(DBGPORT_R11G), .Y(DBG_ADDR722_1)
         );
    zivb U377 ( .A(ADI[9]), .Y(n1081) );
    zmux21lb U378 ( .A(n1072), .B(n1082), .S(DBGPORT_R11G), .Y(DBG_ADDR722_0)
         );
    zivb U379 ( .A(ADI[8]), .Y(n1082) );
    zoai21b U380 ( .A(n1031), .B(n1032), .C(n1033), .Y(DBG_DONE215) );
    zan2b U381 ( .A(DBGPORT_R02G), .B(ADI[16]), .Y(n1031) );
    zmux21lb U382 ( .A(n1042), .B(n1075), .S(DBGPORT_R00G), .Y(DBG_WR403) );
    zivb U383 ( .A(ADI[4]), .Y(n1075) );
    zmux21lb U384 ( .A(n1062), .B(n1083), .S(DBGPORT_R10G), .Y(DBG_ENDP760_3)
         );
    zmux21lb U385 ( .A(n1063), .B(n1054), .S(DBGPORT_R10G), .Y(DBG_ENDP760_2)
         );
    zmux21lb U386 ( .A(n1059), .B(n1080), .S(DBGPORT_R01G), .Y(DBG_INUSE252)
         );
    zivb U387 ( .A(ADI[10]), .Y(n1080) );
    zao32b U388 ( .A(PORT_ENDIS), .B(ADI[28]), .C(DBGPORT_R03G), .D(DBG_ENABLE
        ), .E(n1039), .Y(DBG_ENABLE178) );
    zor2b U389 ( .A(ADI[28]), .B(n1058), .Y(n1039) );
    zivb U390 ( .A(DBGPORT_R03G), .Y(n1058) );
    zmux21lb U391 ( .A(n1038), .B(n1074), .S(DBG_COMPL), .Y(PORT_BLOCK_T326)
         );
    zivb U392 ( .A(PORT_BLOCK), .Y(n1074) );
    zor2b U393 ( .A(PORT_SUSPEND), .B(PORT_RESET), .Y(PORT_BLOCK) );
    zmux21lb U394 ( .A(n1061), .B(n1060), .S(DBG_COMPL), .Y(DBG_ERRGD289) );
    zivb U395 ( .A(DBG_XACTERR), .Y(n1060) );
    zmux21lb U396 ( .A(n1065), .B(n1041), .S(DBGPORT_R10G), .Y(DBG_ENDP760_0)
         );
    zivb U397 ( .A(ADI[0]), .Y(n1041) );
    zmux21hb U398 ( .A(DBG_OWNER), .B(ADI[30]), .S(DBGPORT_R03G), .Y(
        DBG_OWNER141) );
    zan2b U399 ( .A(n1034), .B(n1033), .Y(DBG_GO366) );
    zmux21lb U400 ( .A(n1073), .B(n1050), .S(DBGPORT_R00G), .Y(n1034) );
    zivb U401 ( .A(ADI[5]), .Y(n1050) );
    zivb U402 ( .A(DBG_COMPL), .Y(n1033) );
    zmux21lb U403 ( .A(n1064), .B(n1040), .S(DBGPORT_R10G), .Y(DBG_ENDP760_1)
         );
    zivb U404 ( .A(ADI[1]), .Y(n1040) );
    zan3b U405 ( .A(DBG_ENABLE), .B(n1030), .C(DBGPORT_R03G), .Y(DBG_ENABLE_WC
        ) );
    zivb U406 ( .A(ADI[28]), .Y(n1030) );
    zan2b U407 ( .A(n1085), .B(DBG_TOKEN_0), .Y(DBGPORT_PID[0]) );
    zan2b U408 ( .A(n1085), .B(DBG_TOKEN_1), .Y(DBGPORT_PID[1]) );
    zan2b U409 ( .A(n1085), .B(DBG_TOKEN_2), .Y(DBGPORT_PID[2]) );
    zan2b U410 ( .A(n1085), .B(DBG_TOKEN_3), .Y(DBGPORT_PID[3]) );
    zan2b U411 ( .A(n1085), .B(DBG_TOKEN_4), .Y(DBGPORT_PID[4]) );
    zan2b U412 ( .A(n1085), .B(DBG_TOKEN_5), .Y(DBGPORT_PID[5]) );
    zan2b U413 ( .A(n1028), .B(DBG_TOKEN_6), .Y(DBGPORT_PID[6]) );
    zan2b U414 ( .A(n1085), .B(DBG_TOKEN_7), .Y(DBGPORT_PID[7]) );
    zan2b U415 ( .A(n1028), .B(DBG_TXPID_0), .Y(DBGPORT_PID[8]) );
    zan2b U416 ( .A(n1028), .B(DBG_TXPID_1), .Y(DBGPORT_PID[9]) );
    zan2b U417 ( .A(n1085), .B(DBG_TXPID_2), .Y(DBGPORT_PID[10]) );
    zan2b U418 ( .A(n1085), .B(DBG_TXPID_3), .Y(DBGPORT_PID[11]) );
    zan2b U419 ( .A(n1085), .B(DBG_TXPID_4), .Y(DBGPORT_PID[12]) );
    zan2b U420 ( .A(n1085), .B(DBG_TXPID_5), .Y(DBGPORT_PID[13]) );
    zan2b U421 ( .A(n1028), .B(DBG_TXPID_6), .Y(DBGPORT_PID[14]) );
    zan2b U422 ( .A(n1028), .B(DBG_TXPID_7), .Y(DBGPORT_PID[15]) );
    zan2b U423 ( .A(n1085), .B(DBG_RCVPID_0), .Y(DBGPORT_PID[16]) );
    zan2b U424 ( .A(n1028), .B(DBG_RCVPID_1), .Y(DBGPORT_PID[17]) );
    zan2b U425 ( .A(n1028), .B(DBG_LENGTH_0), .Y(DBGPORT_SC[0]) );
    zan2b U426 ( .A(n1028), .B(DBG_LENGTH_1), .Y(DBGPORT_SC[1]) );
    zan2b U427 ( .A(n1028), .B(DBG_LENGTH_2), .Y(DBGPORT_SC[2]) );
    zan2b U428 ( .A(n1028), .B(DBG_LENGTH_3), .Y(DBGPORT_SC[3]) );
    zan2b U429 ( .A(n1028), .B(DBG_WR), .Y(DBGPORT_SC[4]) );
    zan2b U430 ( .A(DBG_GO), .B(n1028), .Y(DBGPORT_SC[5]) );
    zan2b U431 ( .A(n1028), .B(DBG_ERRGD), .Y(DBGPORT_SC[6]) );
    zan3b U432 ( .A(DBG_XACTERR), .B(n1038), .C(n1084), .Y(DBGPORT_SC[7]) );
    zan3b U433 ( .A(DBG_XACTERR), .B(PORT_BLOCK_T), .C(n1084), .Y(DBGPORT_SC
        [8]) );
    zan2b U434 ( .A(n1028), .B(DBG_INUSE), .Y(DBGPORT_SC[10]) );
    zan2b U435 ( .A(n1028), .B(DBG_DONE), .Y(DBGPORT_SC[16]) );
    zan2b U436 ( .A(n1085), .B(DBG_ENABLE), .Y(DBGPORT_SC[28]) );
    zan2b U437 ( .A(n1085), .B(DBG_OWNER), .Y(DBGPORT_SC[30]) );
    zdffqrb DBG_LENGTH_reg_3 ( .CK(PCICLK_FREE), .D(DBG_LENGTH484_3), .R(n1086
        ), .Q(DBG_LENGTH_3) );
    zdffqrb DBG_LENGTH_reg_2 ( .CK(PCICLK_FREE), .D(DBG_LENGTH484_2), .R(n1087
        ), .Q(DBG_LENGTH_2) );
    zdffqrb DBG_LENGTH_reg_1 ( .CK(PCICLK_FREE), .D(DBG_LENGTH484_1), .R(n1088
        ), .Q(DBG_LENGTH_1) );
    zdffqrb DBG_LENGTH_reg_0 ( .CK(PCICLK_FREE), .D(DBG_LENGTH484_0), .R(n1089
        ), .Q(DBG_LENGTH_0) );
    zdffqrb DBG_RCVPID_reg_7 ( .CK(PCICLK_FREE), .D(DBG_RCVPID572_7), .R(n1086
        ), .Q(DBG_RCVPID_7) );
    zdffqrb DBG_RCVPID_reg_6 ( .CK(PCICLK_FREE), .D(DBG_RCVPID572_6), .R(n1087
        ), .Q(DBG_RCVPID_6) );
    zdffqrb DBG_RCVPID_reg_5 ( .CK(PCICLK_FREE), .D(DBG_RCVPID572_5), .R(n1088
        ), .Q(DBG_RCVPID_5) );
    zdffqrb DBG_RCVPID_reg_4 ( .CK(PCICLK_FREE), .D(DBG_RCVPID572_4), .R(n1089
        ), .Q(DBG_RCVPID_4) );
    zdffqrb DBG_RCVPID_reg_3 ( .CK(PCICLK_FREE), .D(DBG_RCVPID572_3), .R(n1086
        ), .Q(DBG_RCVPID_3) );
    zdffqrb DBG_RCVPID_reg_2 ( .CK(PCICLK_FREE), .D(DBG_RCVPID572_2), .R(n1087
        ), .Q(DBG_RCVPID_2) );
    zdffqrb DBG_RCVPID_reg_1 ( .CK(PCICLK_FREE), .D(DBG_RCVPID572_1), .R(n1088
        ), .Q(DBG_RCVPID_1) );
    zdffqrb DBG_RCVPID_reg_0 ( .CK(PCICLK_FREE), .D(DBG_RCVPID572_0), .R(n1089
        ), .Q(DBG_RCVPID_0) );
    zdffqrb DBG_TXPID_reg_7 ( .CK(PCICLK), .D(DBG_TXPID610_7), .R(n1086), .Q(
        DBG_TXPID_7) );
    zdffqrb DBG_TXPID_reg_6 ( .CK(PCICLK), .D(DBG_TXPID610_6), .R(n1087), .Q(
        DBG_TXPID_6) );
    zivb U438 ( .A(DBG_TXPID_6), .Y(n1043) );
    zdffqrb DBG_TXPID_reg_5 ( .CK(PCICLK), .D(DBG_TXPID610_5), .R(n1088), .Q(
        DBG_TXPID_5) );
    zivb U439 ( .A(DBG_TXPID_5), .Y(n1044) );
    zdffqrb DBG_TXPID_reg_4 ( .CK(PCICLK), .D(DBG_TXPID610_4), .R(n1089), .Q(
        DBG_TXPID_4) );
    zivb U440 ( .A(DBG_TXPID_4), .Y(n1045) );
    zdffqrb DBG_TXPID_reg_3 ( .CK(PCICLK), .D(DBG_TXPID610_3), .R(n1086), .Q(
        DBG_TXPID_3) );
    zivb U441 ( .A(DBG_TXPID_3), .Y(n1046) );
    zdffqrb DBG_TXPID_reg_2 ( .CK(PCICLK), .D(DBG_TXPID610_2), .R(n1087), .Q(
        DBG_TXPID_2) );
    zivb U442 ( .A(DBG_TXPID_2), .Y(n1047) );
    zdffqrb DBG_TXPID_reg_1 ( .CK(PCICLK), .D(DBG_TXPID610_1), .R(n1088), .Q(
        DBG_TXPID_1) );
    zivb U443 ( .A(DBG_TXPID_1), .Y(n1048) );
    zdffqrb DBG_TXPID_reg_0 ( .CK(PCICLK), .D(DBG_TXPID610_0), .R(n1089), .Q(
        DBG_TXPID_0) );
    zivb U444 ( .A(DBG_TXPID_0), .Y(n1049) );
    zdffqrb DBG_TOKEN_reg_7 ( .CK(PCICLK), .D(DBG_TOKEN648_7), .R(n1086), .Q(
        DBG_TOKEN_7) );
    zdffqrb DBG_TOKEN_reg_6 ( .CK(PCICLK), .D(DBG_TOKEN648_6), .R(n1087), .Q(
        DBG_TOKEN_6) );
    zdffqrb DBG_TOKEN_reg_5 ( .CK(PCICLK), .D(DBG_TOKEN648_5), .R(n1088), .Q(
        DBG_TOKEN_5) );
    zivb U445 ( .A(DBG_TOKEN_5), .Y(n1051) );
    zdffqrb DBG_TOKEN_reg_4 ( .CK(PCICLK), .D(DBG_TOKEN648_4), .R(n1089), .Q(
        DBG_TOKEN_4) );
    zivb U446 ( .A(DBG_TOKEN_4), .Y(n1052) );
    zdffqrb DBG_TOKEN_reg_3 ( .CK(PCICLK), .D(DBG_TOKEN648_3), .R(n1086), .Q(
        DBG_TOKEN_3) );
    zivb U447 ( .A(DBG_TOKEN_3), .Y(n1053) );
    zdffqrb DBG_TOKEN_reg_2 ( .CK(PCICLK), .D(DBG_TOKEN648_2), .R(n1087), .Q(
        DBG_TOKEN_2) );
    zivb U448 ( .A(DBG_TOKEN_2), .Y(n1055) );
    zdffqrb DBG_TOKEN_reg_1 ( .CK(PCICLK), .D(DBG_TOKEN648_1), .R(n1088), .Q(
        DBG_TOKEN_1) );
    zivb U449 ( .A(DBG_TOKEN_1), .Y(n1056) );
    zdffqrb DBG_TOKEN_reg_0 ( .CK(PCICLK), .D(DBG_TOKEN648_0), .R(n1089), .Q(
        DBG_TOKEN_0) );
    zivb U450 ( .A(DBG_TOKEN_0), .Y(n1057) );
    zdffqsb DBG_ADDR_reg_6 ( .CK(PCICLK), .D(DBG_ADDR722_6), .S(n1086), .Q(
        DBG_ADDR_6) );
    zivb U451 ( .A(DBG_ADDR_6), .Y(n1066) );
    zdffqsb DBG_ADDR_reg_5 ( .CK(PCICLK), .D(DBG_ADDR722_5), .S(n1087), .Q(
        DBG_ADDR_5) );
    zivb U452 ( .A(DBG_ADDR_5), .Y(n1067) );
    zdffqsb DBG_ADDR_reg_4 ( .CK(PCICLK), .D(DBG_ADDR722_4), .S(n1088), .Q(
        DBG_ADDR_4) );
    zivb U453 ( .A(DBG_ADDR_4), .Y(n1068) );
    zdffqsb DBG_ADDR_reg_3 ( .CK(PCICLK), .D(DBG_ADDR722_3), .S(n1086), .Q(
        DBG_ADDR_3) );
    zivb U454 ( .A(DBG_ADDR_3), .Y(n1069) );
    zdffqsb DBG_ADDR_reg_2 ( .CK(PCICLK), .D(DBG_ADDR722_2), .S(n1087), .Q(
        DBG_ADDR_2) );
    zivb U455 ( .A(DBG_ADDR_2), .Y(n1070) );
    zdffqsb DBG_ADDR_reg_1 ( .CK(PCICLK), .D(DBG_ADDR722_1), .S(n1088), .Q(
        DBG_ADDR_1) );
    zivb U456 ( .A(DBG_ADDR_1), .Y(n1071) );
    zdffqsb DBG_ADDR_reg_0 ( .CK(PCICLK), .D(DBG_ADDR722_0), .S(n1089), .Q(
        DBG_ADDR_0) );
    zivb U457 ( .A(DBG_ADDR_0), .Y(n1072) );
    zdffqrb DBG_DONE_reg ( .CK(PCICLK_FREE), .D(DBG_DONE215), .R(n1086), .Q(
        DBG_DONE) );
    zivb U458 ( .A(DBG_DONE), .Y(n1032) );
    zdffqrb DBG_WR_reg ( .CK(PCICLK), .D(DBG_WR403), .R(n1087), .Q(DBG_WR) );
    zivb U459 ( .A(DBG_WR), .Y(n1042) );
    zdffqrb DBG_ENDP_reg_3 ( .CK(PCICLK), .D(DBG_ENDP760_3), .R(n1088), .Q(
        DBG_ENDP_3) );
    zivb U460 ( .A(DBG_ENDP_3), .Y(n1062) );
    zdffqrb DBG_ENDP_reg_2 ( .CK(PCICLK), .D(DBG_ENDP760_2), .R(n1089), .Q(
        DBG_ENDP_2) );
    zivb U461 ( .A(DBG_ENDP_2), .Y(n1063) );
    zdffqrb DBG_INUSE_reg ( .CK(PCICLK), .D(DBG_INUSE252), .R(n1086), .Q(
        DBG_INUSE) );
    zivb U462 ( .A(DBG_INUSE), .Y(n1059) );
    zdffqrb DBG_ENABLE_reg ( .CK(PCICLK), .D(DBG_ENABLE178), .R(n1087), .Q(
        DBG_ENABLE) );
    zdffqrb PORT_BLOCK_T_reg ( .CK(PCICLK_FREE), .D(PORT_BLOCK_T326), .R(n1088
        ), .Q(PORT_BLOCK_T) );
    zivb U463 ( .A(PORT_BLOCK_T), .Y(n1038) );
    zdffqrb DBG_ERRGD_reg ( .CK(PCICLK_FREE), .D(DBG_ERRGD289), .R(n1089), .Q(
        DBG_ERRGD) );
    zivb U464 ( .A(DBG_ERRGD), .Y(n1061) );
    zdffqsb DBG_ENDP_reg_0 ( .CK(PCICLK), .D(DBG_ENDP760_0), .S(n1086), .Q(
        DBG_ENDP_0) );
    zivb U465 ( .A(DBG_ENDP_0), .Y(n1065) );
    zdffqrb DBG_OWNER_reg ( .CK(PCICLK), .D(DBG_OWNER141), .R(n1086), .Q(
        DBG_OWNER) );
    zdffqrb DBG_GO_reg ( .CK(PCICLK_FREE), .D(DBG_GO366), .R(n1087), .Q(DBG_GO
        ) );
    zivb U466 ( .A(DBG_GO), .Y(n1073) );
    zdffqrb DBG_ENDP_reg_1 ( .CK(PCICLK), .D(DBG_ENDP760_1), .R(n1088), .Q(
        DBG_ENDP_1) );
    zivb U467 ( .A(DBG_ENDP_1), .Y(n1064) );
    znr3b U468 ( .A(DBGPORT_R00G), .B(DBG_WR), .C(n1033), .Y(n1023) );
    zaoi21b U469 ( .A(DBG_COMPL), .B(n1042), .C(DBGPORT_R00G), .Y(n1024) );
    znr2b U470 ( .A(a425), .B(n1041), .Y(n1025) );
    znr2b U471 ( .A(a425), .B(n1040), .Y(n1026) );
    zivb U472 ( .A(ADI[3]), .Y(n1083) );
    zivb U473 ( .A(ADI[2]), .Y(n1054) );
    ziv11b U474 ( .A(EN_DBG_PORT), .Y(n1027), .Z(n1028) );
    zan2b U475 ( .A(n1085), .B(DBG_ADDR_4), .Y(DBGPORT_ADDR[12]) );
    zan2b U476 ( .A(n1084), .B(DBG_ADDR_3), .Y(DBGPORT_ADDR[11]) );
    zan2b U477 ( .A(n1084), .B(DBG_ENDP_2), .Y(DBGPORT_ADDR[2]) );
    zan2b U478 ( .A(n1028), .B(DBG_RCVPID_4), .Y(DBGPORT_PID[20]) );
    zan2b U479 ( .A(n1084), .B(DBG_ENDP_0), .Y(DBGPORT_ADDR[0]) );
    zan2b U480 ( .A(n1084), .B(DBG_RCVPID_6), .Y(DBGPORT_PID[22]) );
    zan2b U481 ( .A(n1084), .B(DBG_RCVPID_2), .Y(DBGPORT_PID[18]) );
    zan2b U482 ( .A(n1084), .B(DBG_ADDR_2), .Y(DBGPORT_ADDR[10]) );
    zan2b U483 ( .A(n1084), .B(DBG_RCVPID_3), .Y(DBGPORT_PID[19]) );
    zan2b U484 ( .A(n1084), .B(DBG_ADDR_5), .Y(DBGPORT_ADDR[13]) );
    zan2b U485 ( .A(n1084), .B(DBG_RCVPID_7), .Y(DBGPORT_PID[23]) );
    zan2b U486 ( .A(n1085), .B(DBG_RCVPID_5), .Y(DBGPORT_PID[21]) );
    zan2b U487 ( .A(n1084), .B(DBG_ENDP_3), .Y(DBGPORT_ADDR[3]) );
    zan2b U488 ( .A(n1084), .B(DBG_ENDP_1), .Y(DBGPORT_ADDR[1]) );
    zan2b U489 ( .A(n1084), .B(DBG_ADDR_0), .Y(DBGPORT_ADDR[8]) );
    zan2b U490 ( .A(n1084), .B(DBG_ADDR_6), .Y(DBGPORT_ADDR[14]) );
    zan2b U491 ( .A(n1084), .B(DBG_ADDR_1), .Y(DBGPORT_ADDR[9]) );
    zivb U492 ( .A(n1027), .Y(n1084) );
    zivb U493 ( .A(n1027), .Y(n1085) );
    zao222b U494 ( .A(DBG_RXBCNT[0]), .B(n1023), .C(DBG_LENGTH_0), .D(n1024), 
        .E(n1025), .F(DBGPORT_R00G), .Y(DBG_LENGTH484_0) );
    zao222b U495 ( .A(DBG_RXBCNT[1]), .B(n1023), .C(DBG_LENGTH_1), .D(n1024), 
        .E(n1026), .F(DBGPORT_R00G), .Y(DBG_LENGTH484_1) );
    zao222b U496 ( .A(DBG_LENGTH_2), .B(n1024), .C(DBG_RXBCNT[2]), .D(n1023), 
        .E(n1035), .F(n1036), .Y(DBG_LENGTH484_2) );
    zao222b U497 ( .A(n1024), .B(DBG_LENGTH_3), .C(n1023), .D(DBG_RXBCNT[3]), 
        .E(DBGPORT_R00G), .F(n1037), .Y(DBG_LENGTH484_3) );
    zbfh U498 ( .A(CMDRST_), .Y(n1086) );
    zbfh U499 ( .A(CMDRST_), .Y(n1087) );
    zbfh U500 ( .A(CMDRST_), .Y(n1088) );
    zbfh U501 ( .A(CMDRST_), .Y(n1089) );
endmodule


// Verilog netlist generated by Chris Lai, 01/17/2000 (13:42:16)

module HS_PCIS (PSADO, FLBASE, CACHLN, ULRDY, UHIT, WR_FRNUM, USBINT, USBEI, 
	HCHALT, USMIO, MAXP, ConfigFlag, FGR, EGSM, GRESET, HCRESET, RUN, 
	UINTOE_, PCI1WAIT, FCFG, PM_EN, HCISPEC_, PAROPT, BABOPT, SUSPORT1, 
	PORTRST1, RESMPRT1, ENPORT1, SUSPORT2, PORTRST2, RESMPRT2, ENPORT2, 
	FB2BKEN, SERREN, RSTEP, RPTYERR, MWRMEN, CAHCFG_, BMASTREN, RDYACK, 
	FRAME0, FRAME4, SOFMOD, REDUCE, /*UDIS1, UDIS2, UENPLL1, UENPLL2, UPD1, 
	UPD2, UTSE01, UTSE02, UTXD1, UTXD2, UTXE1, UTXE2, ULS, UCLK48, URST_, 
	TESTMIA,*/ UIRQSEL3, UIRQSEL2, UIRQSEL1, UIRQSEL0, TESTCNT, ENOCPY, 
	DISEOP, DISPRST, DISSTUFF, /*MIAT,*/ ADI, SERRS, PERRS, MABORTS, TABORTR, 
	CBE3I_, CBE2I_, CBE1I_, CBE0I_, TRDYI_, IRDYI_, FRAMEI_, PMSTR, 
	ERRINT, FRNUM, /*CONN1, CONN2, CONNCHG1, CONNCHG2, CLK_LS,
	ENCHG1, ENCHG2, SDP1, SDP2, SDN1, SDN2, LSDEV1, LSDEV2, RESMDET1, 
	RESMDET2, FGREND, SUSACK1, RESMEND1, ENABLE1, SUSACK2, RESMEND2, 
	ENABLE2, USBRSM, OC1I_, OC0I_, HCHALT_S,*/ HSERR_S, PCIERR_S, ERRINT_S, 
	USBINT_S, FATALINT, RUN_C, CLRHCRST, UADS, /*UCFGCYC,*/ MAC_EOT,
	EHCI_IDLE, PCICLK, PCICLK_FREE, PCIS_ACT, FRNUM_PCLK_LATCH_66,
	HRST_, OCUPY_SEL, DISTXDLY, DISPFUNDRN, ENTXDLY_1, ENTXDLY_2, 
	ENTXDLY_3, SELEOF, DISTXDLY2, DISFFCRC0, DISFFCRC1, DISPFIFO, 
	DISPFIFO2, DISRXZERO, ENBMUSMRST, /*ENLONGPRESOF, DISFFCRC2, DISFFCRC3,
	XUCBE3I_, XUCBE2I_, XUCBE1I_, XUCBE0I_,*/ DEVSELI_, DEVSELO_,
	TRDYO_, TRDYOE_, IDSELI, FUNCSEL, TADOE, TDATA, STOPO_, TPAROE_, LCMD0,
	DISPSTUFF, //DISPLATSOF,		// by Chris Lai, 7/14/2000
	LIGHTRST, ASYNC_EN, PERIOD_EN, ASYNC_ACT, PERIOD_ACT, FRLSTSIZE,
	WR_ASYNCADDR, ASYNCLISTADDR, RECLAMATION, ROLLOVER_S, INTTHRESHOLD,
	/*IOCSPDINT, USBERRINT,*/ USBINT_EN, ERRINT_EN, INTDOORBELL, INTASYNC_EN,
	INTASYNC_S, INTASYNC, ASYNCINT, SLQUEUEADDR, SWDBG, SLAVEMODE,
	SLAVE_ACT, SL_ERROFFSET, CRCERR, PIDERR, SL_DATA_PIDERR,
	SL_ET_ERR, SL_SE_ERR, SL_PCIERR, SL_ACK_ERR, SLAVE_ERR,
	BIST_RUN, BIST_RUN_C, BIST_ERR_S, DIS_BURST,
	TMOUT_PARM, ENISOHANDCHK, DISCHKEOPERR,
	PORTSC1, PORTSC2, PORTSC3, PORTSC4, PORTSC5, PORTSC6, PORTSC7, PORTSC8,
	CFG_CS, PORTCHG_S,

	RxDataOut_A, SquelchOut_A, DisconnectOut_A, TERM_ON_A,
        RxDataOut_B, SquelchOut_B, DisconnectOut_B, TERM_ON_B,
        RxDataOut_C, SquelchOut_C, DisconnectOut_C, TERM_ON_C,
        RxDataOut_D, SquelchOut_D, DisconnectOut_D, TERM_ON_D,
        RxDataOut_E, SquelchOut_E, DisconnectOut_E, TERM_ON_E,
        RxDataOut_F, SquelchOut_F, DisconnectOut_F, TERM_ON_F,
        RxDataOut_G, SquelchOut_G, DisconnectOut_G, TERM_ON_G,
        RxDataOut_H, SquelchOut_H, DisconnectOut_H, TERM_ON_H,

	DIS_TERM_ON_A, DIS_TERM_ON_B, DIS_TERM_ON_C, DIS_TERM_ON_D,
	DIS_TERM_ON_E, DIS_TERM_ON_F, DIS_TERM_ON_G, DIS_TERM_ON_H,
	PSC_CBE2_A, PSC_CBE1_A, PSC_CBE0_A,
        PSC_CBE2_B, PSC_CBE1_B, PSC_CBE0_B,
        PSC_CBE2_C, PSC_CBE1_C, PSC_CBE0_C,
        PSC_CBE2_D, PSC_CBE1_D, PSC_CBE0_D,
        PSC_CBE2_E, PSC_CBE1_E, PSC_CBE0_E,
        PSC_CBE2_F, PSC_CBE1_F, PSC_CBE0_F,
        PSC_CBE2_G, PSC_CBE1_G, PSC_CBE0_G,
        PSC_CBE2_H, PSC_CBE1_H, PSC_CBE0_H,
	R61G, R62G, R63G, R84G, R85G,
	FLADJ5, FLADJ4, FLADJ3, FLADJ2, FLADJ1, FLADJ0,
	PORTWAKECAP8, PORTWAKECAP7, PORTWAKECAP6, PORTWAKECAP5,
	PORTWAKECAP4, PORTWAKECAP3, PORTWAKECAP2, PORTWAKECAP1, PORTWAKECAP0,
	PWR_STATE1, PWR_STATE0, PME_EN, PME_STS, E_PME_EN, PWR_STATE_D0,
        ADS_PRE, LADO,   // by Chris Lai, 1/9/2001
	// USB PHY option bits
	CP0, CP1, SOF_DISCONN_CHK, TEST_FORCE_ENABLE,
        CTRL_A, CTRL_B, CTRL_C, CTRL_D, CTRL_E, CTRL_F, CTRL_G, CTRL_H,
        tst_buferr, loopback, tstmod, rx_block_dis,
        FastLock, LockSpd, TrkSpd, FastStart, RxDataDly, autochk, RDOUT_Enb,
        LBack_Enb, FAST_RST, TMODE, BypassDiv4, UTM_CHKERR,
	sync_fast, sync_jend, SQSET,
	TEST_EYE_EN, FORCE_CRCERR, DIS_NARROW_SOF,
	SetPowner_Dis, PdPHY_Dis, HsEnFB_Dis, ATPG_ENI,
	//FOUNDRYID7, FOUNDRYID6, FOUNDRYID5, FOUNDRYID4,
	//FOUNDRYID3, FOUNDRYID2, FOUNDRYID1, FOUNDRYID0,
	/*EEPHASE, EECFGW0, EECFGW1, EEADO, EECBE,
	EEPA7I, EEPA6I, EEPA5I, EEPA4I, EEPA3I, EEPA2I,
	EECS, EESK, EEDI, EEDO,*/ EN_EHCI, DISPDRCV, CLKOFF_EN, TXTMOUT_EN,
	TXDELAY_EN, TXDELAY_PARM, TURN_PARM, EN_CHKTOGCRC, EN_UTM_RESET,
	EN_REF_RVLD, EN_UTM_SPDUP,
	ENUSB1, ENUSB2, ENUSB3, ENUSB4,
	TRDYOED_, UTM_RUN, SLEEPTIME_SEL,
	BIST_PATTERN, SRAM_WR, SRAM_RUN, SRAM_ADDR, SRAM_SEL,
        SRAM_RDATA1, SRAM_RDATA2, SRAM_RDATA3, SRAM_RDATA4,
	DBGPORT_R08G, DBGPORT_R09G, DBGPORT_R0AG, DBGPORT_R0BG,
	DBGPORT_R0CG, DBGPORT_R0DG, DBGPORT_R0EG, DBGPORT_R0FG,
	EN_DBG_PORT, DBGPORT_SC, DBGPORT_PID, DBGPORT_ADDR,
	DBGPORT_BUF1, DBGPORT_BUF2, DBG_COMPL, DBG_XACTERR,
	DBG_RXBCNT, DBG_RXPID, DBG_ENABLE_WC );
output	DBGPORT_R08G, DBGPORT_R09G, DBGPORT_R0AG, DBGPORT_R0BG,
        DBGPORT_R0CG, DBGPORT_R0DG, DBGPORT_R0EG, DBGPORT_R0FG,
	EN_DBG_PORT, DBG_ENABLE_WC;
output	[31:0]	DBGPORT_SC, DBGPORT_PID, DBGPORT_ADDR;
input	[31:0]	DBGPORT_BUF1, DBGPORT_BUF2;
input	DBG_COMPL, DBG_XACTERR;
input	[3:0]	DBG_RXBCNT;
input	[7:0]	DBG_RXPID;
input	FRNUM_PCLK_LATCH_66;
output	sync_fast, sync_jend;
output	[1:0]	SQSET;
output  [31:0]  BIST_PATTERN;
output  [8:0]   SRAM_ADDR;
output  [1:0]   SRAM_SEL;
output          SRAM_WR, SRAM_RUN;
input   [31:0]  SRAM_RDATA1, SRAM_RDATA2, SRAM_RDATA3, SRAM_RDATA4;
output	TRDYOED_, UTM_RUN, SLEEPTIME_SEL;
input	ENUSB1, ENUSB2, ENUSB3, ENUSB4;
output	EN_CHKTOGCRC, EN_UTM_RESET, EN_REF_RVLD, EN_UTM_SPDUP;
output	/*EEPHASE, EECFGW0, EECFGW1, EECS, EESK, EEDI,*/ UADS, TXTMOUT_EN;
output	/*EEPA7I, EEPA6I, EEPA5I, EEPA4I, EEPA3I, EEPA2I,*/ DISPDRCV, CLKOFF_EN;
input	/*EEDO,*/ EN_EHCI;
//output	[31:0]	EEADO;
//output	[3:0]	EECBE;
output  CP0, CP1, SOF_DISCONN_CHK, loopback, tstmod, rx_block_dis, tst_buferr,
        RDOUT_Enb, FastLock, LBack_Enb, FAST_RST, TMODE, FastStart, BypassDiv4;
output	autochk, SetPowner_Dis, PdPHY_Dis, HsEnFB_Dis;
output  [3:0]   CTRL_A, CTRL_B, CTRL_C, CTRL_D, CTRL_E, CTRL_F, CTRL_G, CTRL_H;
output  [2:0]   RxDataDly;
output  [1:0]   LockSpd, TrkSpd;
output	[7:0]	TMOUT_PARM, TXDELAY_PARM;
output	[3:0]	TURN_PARM;
output	TXDELAY_EN;
output	ENISOHANDCHK, DISCHKEOPERR;
output	ADS_PRE;
output	[31:0]	LADO;
output	R61G, R62G, R63G, R84G, R85G;
input	FLADJ5, FLADJ4, FLADJ3, FLADJ2, FLADJ1, FLADJ0,
	PORTWAKECAP8, PORTWAKECAP7, PORTWAKECAP6, PORTWAKECAP5,
	PORTWAKECAP4, PORTWAKECAP3, PORTWAKECAP2, PORTWAKECAP1, PORTWAKECAP0,
	PWR_STATE1, PWR_STATE0, PME_EN, PME_STS, E_PME_EN, PWR_STATE_D0;
input	BIST_RUN_C, BIST_ERR_S, UTM_CHKERR;
output	BIST_RUN, DIS_BURST, TEST_EYE_EN, FORCE_CRCERR, DIS_NARROW_SOF;
input	CRCERR, PIDERR, SL_DATA_PIDERR, SL_ET_ERR, SL_SE_ERR, SL_ACK_ERR;
input	SL_PCIERR, SLAVE_ERR;
output	[31:0]	SLQUEUEADDR;
output	SWDBG, SLAVEMODE;
input	SLAVE_ACT;
input	[7:0]	SL_ERROFFSET;
input	INTASYNC_S, ASYNCINT;
output	USBINT_EN, ERRINT_EN, INTASYNC_EN, INTDOORBELL, INTASYNC;
//input	IOCSPDINT, USBERRINT;
output	[7:0]	INTTHRESHOLD;
output	LIGHTRST, ASYNC_EN, PERIOD_EN, WR_ASYNCADDR;
input	ASYNC_ACT, PERIOD_ACT, RECLAMATION, ROLLOVER_S, EHCI_IDLE;
output	[1:0]	FRLSTSIZE;
input	[31:0]	ASYNCLISTADDR;
output	DISPSTUFF; //DISFFCRC3, DISPLATSOF;	// by Chris Lai, 7/14/2000
output	TADOE, TDATA, STOPO_, TPAROE_, LCMD0;
input	DEVSELI_, IDSELI;//, FUNCSEL;
input	[2:0] FUNCSEL;
output	DEVSELO_, TRDYO_, TRDYOE_;
output	[31:0]	PSADO;
output	[31:12]	FLBASE;
output	[7:0]	CACHLN;
output	ULRDY, UHIT, WR_FRNUM, USBINT, USBEI, HCHALT, USMIO, MAXP;
output	FGR, EGSM, GRESET, HCRESET, RUN, UINTOE_, PCI1WAIT, FCFG, PM_EN;
output	HCISPEC_, PAROPT, BABOPT, SUSPORT1, PORTRST1, RESMPRT1, ENPORT1;
output	SUSPORT2, PORTRST2, RESMPRT2, ENPORT2, FB2BKEN, SERREN, RSTEP;
output	RPTYERR, MWRMEN, CAHCFG_, BMASTREN, RDYACK, FRAME0, FRAME4;
output	[7:0]	SOFMOD;
//output	REDUCE, UDIS1, UDIS2, UENPLL1, UENPLL2, UPD1, UPD2, UTSE01, UTSE02;
//output	UTXD1, UTXD2, UTXE1, UTXE2, ULS, UCLK48, URST_, TESTMIA, UIRQSEL3;
output	REDUCE, UIRQSEL3;
output	UIRQSEL2, UIRQSEL1, UIRQSEL0, TESTCNT, ENOCPY, DISEOP, DISPRST;
output	DISSTUFF;
//input	[31:1]	MIAT;
input	[31:0]	ADI;
input	SERRS, PERRS, MABORTS, TABORTR, CBE3I_, CBE2I_, CBE1I_, CBE0I_;
input	TRDYI_, IRDYI_, FRAMEI_, PMSTR;//, IOCINT, SPDINT;//
output	ERRINT;
input	[13:0]	FRNUM;
/*
input	CONN1, CONN2, CONNCHG1, CONNCHG2, ENCHG1, ENCHG2, SDP1, SDP2, SDN1;
input	SDN2, LSDEV1, LSDEV2, RESMDET1, RESMDET2, FGREND, SUSACK1, RESMEND1;
input	ENABLE1, SUSACK2, RESMEND2, ENABLE2, USBRSM, OC1I_, OC0I_;*/
input	HSERR_S, PCIERR_S, ERRINT_S, USBINT_S, FATALINT, RUN_C, CLRHCRST;
input	/*UADS, UCFGCYC,*/ MAC_EOT, PCICLK, PCICLK_FREE, HRST_;//, HCHALT_S, CLK_LS;
output	PCIS_ACT;
output	[1:0]	OCUPY_SEL;
output	DISTXDLY, DISPFUNDRN, ENTXDLY_1, ENTXDLY_2, ENTXDLY_3, SELEOF;
output	DISTXDLY2, DISFFCRC0, DISFFCRC1, DISPFIFO, DISPFIFO2, DISRXZERO;
output	ENBMUSMRST;//, ENLONGPRESOF;//, DISFFCRC2;
input	ConfigFlag;
input	[31:0]	PORTSC1, PORTSC2, PORTSC3, PORTSC4, PORTSC5, PORTSC6,
		PORTSC7, PORTSC8;
output	CFG_CS;
output	PSC_CBE2_A, PSC_CBE1_A, PSC_CBE0_A,
        PSC_CBE2_B, PSC_CBE1_B, PSC_CBE0_B,
        PSC_CBE2_C, PSC_CBE1_C, PSC_CBE0_C,
        PSC_CBE2_D, PSC_CBE1_D, PSC_CBE0_D,
        PSC_CBE2_E, PSC_CBE1_E, PSC_CBE0_E,
        PSC_CBE2_F, PSC_CBE1_F, PSC_CBE0_F,
        PSC_CBE2_G, PSC_CBE1_G, PSC_CBE0_G,
        PSC_CBE2_H, PSC_CBE1_H, PSC_CBE0_H;
input	TEST_FORCE_ENABLE, PORTCHG_S;
input   RxDataOut_A, SquelchOut_A, DisconnectOut_A, TERM_ON_A,
        RxDataOut_B, SquelchOut_B, DisconnectOut_B, TERM_ON_B,
        RxDataOut_C, SquelchOut_C, DisconnectOut_C, TERM_ON_C,
        RxDataOut_D, SquelchOut_D, DisconnectOut_D, TERM_ON_D,
        RxDataOut_E, SquelchOut_E, DisconnectOut_E, TERM_ON_E,
        RxDataOut_F, SquelchOut_F, DisconnectOut_F, TERM_ON_F,
        RxDataOut_G, SquelchOut_G, DisconnectOut_G, TERM_ON_G,
        RxDataOut_H, SquelchOut_H, DisconnectOut_H, TERM_ON_H;
output	DIS_TERM_ON_A, DIS_TERM_ON_B, DIS_TERM_ON_C, DIS_TERM_ON_D,
	DIS_TERM_ON_E, DIS_TERM_ON_F, DIS_TERM_ON_G, DIS_TERM_ON_H;
//input	FOUNDRYID7, FOUNDRYID6, FOUNDRYID5, FOUNDRYID4,
//	FOUNDRYID3, FOUNDRYID2, FOUNDRYID1, FOUNDRYID0;
input	ATPG_ENI;
//input	XUCBE3I_, XUCBE2I_, XUCBE1I_, XUCBE0I_;
/*wire	CFGW, REGW, 
	REGR, REGADS, REGD31, 
	REGD30, REGD29, REGD28, REGD27, REGD26, REGD25, REGD24, REGD23, REGD22, 
	REGD21, REGD20, REGD19, REGD18, REGD17, REGD16, REGD15, REGD14, REGD13, 
	REGD12, REGD11, REGD10, REGD9, REGD8, REGD7, REGD6, REGD5, REGD4, 
	REGD3, REGD2, REGD1, REGD0, CFGD31, CFGD30, CFGD29, CFGD28, CFGD27, 
	CFGD26, CFGD25, CFGD24, CFGD23, CFGD22, CFGD21, CFGD20, CFGD19, CFGD18, 
	CFGD17, CFGD16, CFGD15, CFGD14, CFGD13, CFGD12, CFGD11, CFGD10, CFGD9, 
	CFGD8, CFGD7, CFGD6, CFGD5, CFGD4, CFGD3, CFGD2, CFGD1, CFGD0, IOBA31, 
	IOBA30, IOBA29, IOBA28, IOBA27, IOBA26, IOBA25, IOBA24, IOBA23, IOBA22, 
	IOBA21, IOBA20, IOBA19, IOBA18, IOBA17, IOBA16, IOBA15, IOBA14, IOBA13, 
	IOBA12, IOBA11, IOBA10, IOBA9, IOBA8, 
	VIAPSS, UIRQACT, 
	IOSPACE, DEVS0, MMSPACE, DBGIRQ, UIRQEN, USBSPEC7, USBSPEC6, USBSPEC5, 
	USBSPEC4, USBSPEC3, USBSPEC2, USBSPEC1, USBSPEC0, REVID7, REVID6, 
	REVID5, REVID4, REVID3, REVID2, REVID1, REVID0, MAXLAT7, MAXLAT6, 
	MAXLAT5, MAXLAT4, MAXLAT3, MAXLAT2, MAXLAT1, MAXLAT0, MINGNT7, MINGNT6, 
	MINGNT5, MINGNT4, MINGNT3, MINGNT2, MINGNT1, MINGNT0;*/
wire	[31:0] LADO;
wire	[3:0] LCBE;
/*wire	ADS, LCMD0, PA7I, PA6I, PA5I, PA4I, PA3I, PA2I, THIT, ADRG, TADOE, 
	TERM, TDATA, TRDYO_, STOPO_, DEVSELO_, TRDYOE_, TPAROE_, DEVSELI_, HIT, 
	LRDY, TGWR;*/
wire [31:0] USBLEGCTLSTS, USBLEGSUP;
//wire [5:0]  EEP_ADDR;
//wire [15:0] EEP_RDATA;
//wire [31:0] ULADO, EEADO;
//wire [3:0]  ULCBE, EECBE;
wire VDD = 1'b1;
wire GND = 1'b0;
    ULAD ULAD ( .ADI({ADI[31], ADI[30], ADI[29], ADI[28], ADI[27], ADI[26], 
	ADI[25], ADI[24], ADI[23], ADI[22], ADI[21], ADI[20], ADI[19], ADI[18]
	, ADI[17], ADI[16], ADI[15], ADI[14], ADI[13], ADI[12], ADI[11], 
	ADI[10], ADI[9], ADI[8], ADI[7], ADI[6], ADI[5], ADI[4], ADI[3], 
	ADI[2], ADI[1], ADI[0]}), .CBEI_({CBE3I_, CBE2I_, CBE1I_, CBE0I_}), 
	.ADS_PRE(ADS_PRE), .HRST_(HRST_),.LADO({LADO[31], LADO[30], LADO[29], 
	LADO[28], LADO[27], LADO[26], LADO[25], LADO[24], LADO[23], LADO[22], 
	LADO[21], LADO[20], LADO[19], LADO[18], LADO[17], LADO[16], LADO[15], 
	LADO[14], LADO[13], LADO[12], LADO[11], LADO[10], LADO[9], LADO[8], 
	LADO[7], LADO[6], LADO[5], LADO[4], LADO[3], LADO[2], LADO[1], LADO[0]
	}), .LCBE({LCBE[3], LCBE[2], LCBE[1], LCBE[0]}),
	/*.LADO(ULADO), .LCBE(ULCBE),*/ .PCICLK(PCICLK) );
    HS_INTF HS_INTF ( .PSADO31(PSADO[31]), .PSADO30(PSADO[30]), .PSADO29(PSADO[29]
	), .PSADO28(PSADO[28]), .PSADO27(PSADO[27]), .PSADO26(PSADO[26]), 
	.PSADO25(PSADO[25]), .PSADO24(PSADO[24]), .PSADO23(PSADO[23]), 
	.PSADO22(PSADO[22]), .PSADO21(PSADO[21]), .PSADO20(PSADO[20]), 
	.PSADO19(PSADO[19]), .PSADO18(PSADO[18]), .PSADO17(PSADO[17]), 
	.PSADO16(PSADO[16]), .PSADO15(PSADO[15]), .PSADO14(PSADO[14]), 
	.PSADO13(PSADO[13]), .PSADO12(PSADO[12]), .PSADO11(PSADO[11]), 
	.PSADO10(PSADO[10]), .PSADO9(PSADO[9]), .PSADO8(PSADO[8]), .PSADO7(
	PSADO[7]), .PSADO6(PSADO[6]), .PSADO5(PSADO[5]), .PSADO4(PSADO[4]), 
	.PSADO3(PSADO[3]), .PSADO2(PSADO[2]), .PSADO1(PSADO[1]), .PSADO0(
	PSADO[0]), .UHIT(UHIT),
	.ULRDY(ULRDY), .CFGW(CFGW), .REGW(REGW), .REGR(REGR), .REGADS(
	//.ULRDY(ULRDY), .CFGW(UCFGW), .REGW(REGW), .REGR(REGR), .REGADS(
	REGADS), .RDYACK(RDYACK), 
	.IRDYI_(IRDYI_), 
	.TRDYI_(TRDYI_), /*.FRAMEI_(FRAMEI_),*/.LCMD0(LCMD0), .AD31I(ADI[31]), 
	.AD30I(ADI[30]), .AD29I(ADI[29]), .AD28I(ADI[28]), .AD27I(ADI[27]), 
	.AD26I(ADI[26]), .AD25I(ADI[25]), .AD24I(ADI[24]), .AD23I(ADI[23]), 
	.AD22I(ADI[22]), .AD21I(ADI[21]), .AD20I(ADI[20]), .AD19I(ADI[19]), 
	.AD18I(ADI[18]), .AD17I(ADI[17]), .AD16I(ADI[16]), .AD15I(ADI[15]), 
	.AD14I(ADI[14]), .AD13I(ADI[13]), .AD12I(ADI[12]), .AD11I(ADI[11]), 
	.AD10I(ADI[10]), .AD9I(ADI[9]), .AD8I(ADI[8]), .AD7I(ADI[7]), .AD6I(
	ADI[6]), .AD5I(ADI[5]), .AD4I(ADI[4]), .AD3I(ADI[3]), .AD2I(ADI[2]), 
	.AD1I(ADI[1]), .AD0I(ADI[0]), .REGD31(REGD31), .REGD30(REGD30), 
	.REGD29(REGD29), .REGD28(REGD28), .REGD27(REGD27), .REGD26(REGD26), 
	.REGD25(REGD25), .REGD24(REGD24), .REGD23(REGD23), .REGD22(REGD22), 
	.REGD21(REGD21), .REGD20(REGD20), .REGD19(REGD19), .REGD18(REGD18), 
	.REGD17(REGD17), .REGD16(REGD16), .REGD15(REGD15), .REGD14(REGD14), 
	.REGD13(REGD13), .REGD12(REGD12), .REGD11(REGD11), .REGD10(REGD10), 
	.REGD9(REGD9), .REGD8(REGD8), .REGD7(REGD7), .REGD6(REGD6), .REGD5(
	REGD5), .REGD4(REGD4), .REGD3(REGD3), .REGD2(REGD2), .REGD1(REGD1), 
	.REGD0(REGD0), .CFGD31(CFGD31), .CFGD30(CFGD30), .CFGD29(CFGD29), 
	.CFGD28(CFGD28), .CFGD27(CFGD27), .CFGD26(CFGD26), .CFGD25(CFGD25), 
	.CFGD24(CFGD24), .CFGD23(CFGD23), .CFGD22(CFGD22), .CFGD21(CFGD21), 
	.CFGD20(CFGD20), .CFGD19(CFGD19), .CFGD18(CFGD18), .CFGD17(CFGD17), 
	.CFGD16(CFGD16), .CFGD15(CFGD15), .CFGD14(CFGD14), .CFGD13(CFGD13), 
	.CFGD12(CFGD12), .CFGD11(CFGD11), .CFGD10(CFGD10), .CFGD9(CFGD9), 
	.CFGD8(CFGD8), .CFGD7(CFGD7), .CFGD6(CFGD6), .CFGD5(CFGD5), .CFGD4(
	CFGD4), .CFGD3(CFGD3), .CFGD2(CFGD2), .CFGD1(CFGD1), .CFGD0(CFGD0), 
	.CBE3I_(CBE3I_), .CBE2I_(CBE2I_), .CBE1I_(CBE1I_), .CBE0I_(
	CBE0I_), .IOBA31(IOBA31), .IOBA30(IOBA30), .IOBA29(IOBA29), .IOBA28(
	IOBA28), .IOBA27(IOBA27), .IOBA26(IOBA26), .IOBA25(IOBA25), .IOBA24(
	IOBA24), .IOBA23(IOBA23), .IOBA22(IOBA22), .IOBA21(IOBA21), .IOBA20(
	IOBA20), .IOBA19(IOBA19), .IOBA18(IOBA18), .IOBA17(IOBA17), .IOBA16(
	IOBA16), .IOBA15(IOBA15), .IOBA14(IOBA14), .IOBA13(IOBA13), .IOBA12(
	IOBA12), .IOBA11(IOBA11), .IOBA10(IOBA10), .IOBA9(IOBA9),
	.IOBA8(IOBA8),  //.UIRQACT(UIRQACT), 
	//.UADS(UADS), /*.UCFGCYC(UCFGCYC),*/ .IOSPACE(IOSPACE), .PMSTR(PMSTR), 
	.UADS(UADS), /*.UCFGCYC(UCFGCYC),*/ .IOSPACE(MMSPACE), .PMSTR(PMSTR), 
	.HRST_(HRST_), .PCICLK(PCICLK_FREE), .ADS(ADS), .ADRG(ADRG), .PA7I(PA7I), 
	.PA6I(PA6I), .PA5I(PA5I), .PA4I(PA4I), .PA3I(PA3I), .PA2I(PA2I),
	.FUNCSEL(FUNCSEL), .IDSELI(IDSELI), .EN_EHCI(EN_EHCI) );

// Foundry ID => 03 (TSMC fab.4)
//smux21id        DNTFID0(.Y(FOUNDRYID0),.A(VDD),.B(GND),.S(VDD));
//smux21id        DNTFID1(.Y(FOUNDRYID1),.A(VDD),.B(GND),.S(VDD));
//smux21id        DNTFID2(.Y(FOUNDRYID2),.A(VDD),.B(GND),.S(GND));
//smux21id        DNTFID3(.Y(FOUNDRYID3),.A(VDD),.B(GND),.S(GND));
//smux21id        DNTFID4(.Y(FOUNDRYID4),.A(VDD),.B(GND),.S(GND));
//smux21id        DNTFID5(.Y(FOUNDRYID5),.A(VDD),.B(GND),.S(GND));
//smux21id        DNTFID6(.Y(FOUNDRYID6),.A(VDD),.B(GND),.S(GND));
//smux21id        DNTFID7(.Y(FOUNDRYID7),.A(VDD),.B(GND),.S(GND));

    HS_PCICFG HS_PCICFG ( .CFGD31(CFGD31), .CFGD30(CFGD30), .CFGD29(CFGD29), 
	.CFGD28(CFGD28), .CFGD27(CFGD27), .CFGD26(CFGD26), .CFGD25(CFGD25), 
	.CFGD24(CFGD24), .CFGD23(CFGD23), .CFGD22(CFGD22), .CFGD21(CFGD21), 
	.CFGD20(CFGD20), .CFGD19(CFGD19), .CFGD18(CFGD18), .CFGD17(CFGD17), 
	.CFGD16(CFGD16), .CFGD15(CFGD15), .CFGD14(CFGD14), .CFGD13(CFGD13), 
	.CFGD12(CFGD12), .CFGD11(CFGD11), .CFGD10(CFGD10), .CFGD9(CFGD9), 
	.CFGD8(CFGD8), .CFGD7(CFGD7), .CFGD6(CFGD6), .CFGD5(CFGD5), .CFGD4(
	CFGD4), .CFGD3(CFGD3), .CFGD2(CFGD2), .CFGD1(CFGD1), .CFGD0(CFGD0), 
	.IOBA31(IOBA31), .IOBA30(IOBA30), .IOBA29(IOBA29), .IOBA28(IOBA28), 
	.IOBA27(IOBA27), .IOBA26(IOBA26), .IOBA25(IOBA25), .IOBA24(IOBA24), 
	.IOBA23(IOBA23), .IOBA22(IOBA22), .IOBA21(IOBA21), .IOBA20(IOBA20), 
	.IOBA19(IOBA19), .IOBA18(IOBA18), .IOBA17(IOBA17), .IOBA16(IOBA16), 
	.IOBA15(IOBA15), .IOBA14(IOBA14), .IOBA13(IOBA13), .IOBA12(IOBA12), 
	.IOBA11(IOBA11), .IOBA10(IOBA10), .IOBA9(IOBA9), .IOBA8(IOBA8), 
	.CACHLN7(CACHLN[7]), 
	.CACHLN6(CACHLN[6]), .CACHLN5(CACHLN[5]), .CACHLN4(CACHLN[4]), 
	.CACHLN3(CACHLN[3]), .CACHLN2(CACHLN[2]), .CACHLN1(CACHLN[1]), 
	.CACHLN0(CACHLN[0]), .DEVS0(DEVS0), .FB2BKEN(FB2BKEN), .SERREN(SERREN)
	, .RSTEP(RSTEP), .RPTYERR(RPTYERR), .MWRMEN(MWRMEN), .BMASTREN(
	BMASTREN), .MMSPACE(MMSPACE), .IOSPACE(IOSPACE), .UIRQSEL3(UIRQSEL3), 
	.UIRQSEL2(UIRQSEL2), .UIRQSEL1(UIRQSEL1), .UIRQSEL0(UIRQSEL0), 
	.PCI1WAIT(PCI1WAIT), .FCFG(FCFG), .PM_EN(PM_EN), .HCISPEC_(HCISPEC_), 
	.REDUCE(REDUCE), .PAROPT(PAROPT), .BABOPT(BABOPT), .CAHCFG_(CAHCFG_), 
	.TRAP_OPT(TRAP_OPT), .VIAPSS(VIAPSS), .DBGIRQ(DBGIRQ), /*.UDIS1(UDIS1), 
	.UDIS2(UDIS2), .UENPLL1(UENPLL1), .UENPLL2(UENPLL2), .UPD1(UPD1), 
	.UPD2(UPD2), .UTSE01(UTSE01), .UTSE02(UTSE02), .UTXD1(UTXD1), .UTXD2(
	UTXD2), .UTXE1(UTXE1), .UTXE2(UTXE2), .ULS(ULS), .UCLK48(UCLK48), 
	.URST_(URST_), .TESTMIA(TESTMIA),*/ .ENOCPY(ENOCPY), .DISEOP(DISEOP), 
	.DISPRST(DISPRST), .DISSTUFF(DISSTUFF),
	.TESTCNT(TESTCNT), 
	/*.MIAT31(MIAT[31]), .MIAT30(MIAT[30]), .MIAT29(MIAT[29]), .MIAT28(
	MIAT[28]), .MIAT27(MIAT[27]), .MIAT26(MIAT[26]), .MIAT25(MIAT[25]), 
	.MIAT24(MIAT[24]), .MIAT23(MIAT[23]), .MIAT22(MIAT[22]), .MIAT21(
	MIAT[21]), .MIAT20(MIAT[20]), .MIAT19(MIAT[19]), .MIAT18(MIAT[18]), 
	.MIAT17(MIAT[17]), .MIAT16(MIAT[16]), .MIAT15(MIAT[15]), .MIAT14(
	MIAT[14]), .MIAT13(MIAT[13]), .MIAT12(MIAT[12]), .MIAT11(MIAT[11]), 
	.MIAT10(MIAT[10]), .MIAT09(MIAT[9]), .MIAT08(MIAT[8]), .MIAT07(MIAT[7]
	), .MIAT06(MIAT[6]), .MIAT05(MIAT[5]), .MIAT04(MIAT[4]), .MIAT03(
	MIAT[3]), .MIAT02(MIAT[2]), .MIAT01(MIAT[1]),*/ .AD31I(LADO[31]), 
	.AD30I(LADO[30]), .AD29I(LADO[29]), .AD28I(LADO[28]), .AD27I(LADO[27])
	, .AD26I(LADO[26]), .AD25I(LADO[25]), .AD24I(LADO[24]), .AD23I(
	LADO[23]), .AD22I(LADO[22]), .AD21I(LADO[21]), .AD20I(LADO[20]), 
	.AD19I(LADO[19]), .AD18I(LADO[18]), .AD17I(LADO[17]), .AD16I(LADO[16])
	, .AD15I(LADO[15]), .AD14I(LADO[14]), .AD13I(LADO[13]), .AD12I(
	LADO[12]), .AD11I(LADO[11]), .AD10I(LADO[10]), .AD9I(LADO[9]), .AD8I(
	LADO[8]), .AD7I(LADO[7]), .AD6I(LADO[6]), .AD5I(LADO[5]), .AD4I(
	LADO[4]), .AD3I(LADO[3]), .AD2I(LADO[2]), .AD1I(LADO[1]), .AD0I(
	LADO[0]), .PA7I(PA7I), .PA6I(PA6I), .PA5I(PA5I), .PA4I(PA4I), .PA3I(
	PA3I), .PA2I(PA2I), .CBE3I_(LCBE[3]), .CBE2I_(LCBE[2]), .CBE1I_(
	LCBE[1]), .CBE0I_(LCBE[0]), .CFGW(CFGW),
	/*.USBSPEC7(USBSPEC7), .USBSPEC6(USBSPEC6), .USBSPEC5(USBSPEC5),
	.USBSPEC4(USBSPEC4), .USBSPEC3(USBSPEC3), .USBSPEC2(USBSPEC2),
	.USBSPEC1(USBSPEC1), .USBSPEC0(USBSPEC0),*/
	.REVID7(REVID7), .REVID6(REVID6), .REVID5(REVID5), .REVID4(REVID4),
	.REVID3(REVID3), .REVID2(REVID2), .REVID1(REVID1), .REVID0(REVID0),
	/*.FOUNDRYID0(FOUNDRYID0), .FOUNDRYID1(FOUNDRYID1),
	.FOUNDRYID2(FOUNDRYID2), .FOUNDRYID3(FOUNDRYID3),
	.FOUNDRYID4(FOUNDRYID4), .FOUNDRYID5(FOUNDRYID5),
	.FOUNDRYID6(FOUNDRYID6), .FOUNDRYID7(FOUNDRYID7),*/
	.MAXLAT7(MAXLAT7), .MAXLAT6(MAXLAT6), .MAXLAT5(MAXLAT5),
	.MAXLAT4(MAXLAT4), .MAXLAT3(MAXLAT3), .MAXLAT2(MAXLAT2), 
	.MAXLAT1(MAXLAT1), .MAXLAT0(MAXLAT0), .MINGNT7(MINGNT7), .MINGNT6(
	MINGNT6), .MINGNT5(MINGNT5), .MINGNT4(MINGNT4), .MINGNT3(MINGNT3), 
	.MINGNT2(MINGNT2), .MINGNT1(MINGNT1), .MINGNT0(MINGNT0), 
	.UIRQACT(UIRQACT), .SERRS(SERRS), 
	.MABORTS(MABORTS), .TABORTR(TABORTR),
	.INTR_DIS(INTR_DIS),
	.PCICLK(PCICLK), .PCICLK_FREE(PCICLK_FREE), .HRST_(HRST_), 
	.OCUPY_SEL({OCUPY_SEL[1], OCUPY_SEL[0]}), .DISTXDLY(DISTXDLY), 
	.DISPFUNDRN(DISPFUNDRN), .ENTXDLY_1(ENTXDLY_1), .ENTXDLY_2(ENTXDLY_2)
	, .ENTXDLY_3(ENTXDLY_3), .SELEOF(SELEOF), .DISTXDLY2(DISTXDLY2), 
	.DISFFCRC0(DISFFCRC0), .DISFFCRC1(DISFFCRC1), .DISPFIFO(DISPFIFO), 
	.DISPFIFO2(DISPFIFO2), .DISRXZERO(DISRXZERO), .ENBMUSMRST(ENBMUSMRST)
	, /*.DISFFCRC2(DISFFCRC2), .ENLONGPRESOF(ENLONGPRESOF),*/
	.FUNCSEL(FUNCSEL), /*.DISFFCRC3(DISFFCRC3),*/ .DISPSTUFF(DISPSTUFF),
	//.DISPLATSOF(DISPLATSOF),	// by Chris Lai, 7/14/2000
	.HCHALT(HCHALT), .CMDRST_(CMDRST_), .SWDBG(SWDBG),
	.SLQUEUEADDR(SLQUEUEADDR), .SLAVEMODE(SLAVEMODE),
	.SLAVE_ACT(SLAVE_ACT), .SL_ERROFFSET(SL_ERROFFSET),
	.CRCERR(CRCERR), .PIDERR(PIDERR), .SL_DATA_PIDERR(SL_DATA_PIDERR),
	.SL_ET_ERR(SL_ET_ERR), .SL_SE_ERR(SL_SE_ERR), .SL_PCIERR(SL_PCIERR),
	.SL_ACK_ERR(SL_ACK_ERR), .SLAVE_ERR(SLAVE_ERR),
	.BIST_RUN(BIST_RUN), .BIST_RUN_C(BIST_RUN_C),
	.BIST_ERR_S(BIST_ERR_S), .DIS_BURST(DIS_BURST),
	.TMOUT_PARM(TMOUT_PARM), .ENISOHANDCHK(ENISOHANDCHK),
	.DISCHKEOPERR(DISCHKEOPERR), .EN_CHKTOGCRC(EN_CHKTOGCRC),
	.EN_UTM_RESET(EN_UTM_RESET), .EN_REF_RVLD(EN_REF_RVLD),
	.EN_UTM_SPDUP(EN_UTM_SPDUP),
	.R61G(R61G), .R62G(R62G), .R63G(R63G), .R84G(R84G), .R85G(R85G),
	.FLADJ5(FLADJ5), .FLADJ4(FLADJ4), .FLADJ3(FLADJ3), .FLADJ2(FLADJ2),
	.FLADJ1(FLADJ1), .FLADJ0(FLADJ0), .PORTWAKECAP8(PORTWAKECAP8),
	.PORTWAKECAP7(PORTWAKECAP7), .PORTWAKECAP6(PORTWAKECAP6),
	.PORTWAKECAP5(PORTWAKECAP5), .PORTWAKECAP4(PORTWAKECAP4),
	.PORTWAKECAP3(PORTWAKECAP3), .PORTWAKECAP2(PORTWAKECAP2),
	.PORTWAKECAP1(PORTWAKECAP1), .PORTWAKECAP0(PORTWAKECAP0),
	.PWR_STATE1(PWR_STATE1), .PWR_STATE0(PWR_STATE0),
	.PME_EN(PME_EN), .PME_STS(PME_STS), .E_PME_EN(E_PME_EN),
	.CP0(CP0), .CP1(CP1), .SOF_DISCONN_CHK(SOF_DISCONN_CHK),
	.CTRL_A(CTRL_A), .CTRL_B(CTRL_B), .CTRL_C(CTRL_C), .CTRL_D(CTRL_D),
	.CTRL_E(CTRL_E), .CTRL_F(CTRL_F), .CTRL_G(CTRL_G), .CTRL_H(CTRL_H),
	.loopback(loopback), .tstmod(tstmod), .rx_block_dis(rx_block_dis),
	.FastLock(FastLock), .LockSpd(LockSpd), .TrkSpd(TrkSpd),
	.RxDataDly(RxDataDly), .RDOUT_Enb(RDOUT_Enb), .LBack_Enb(LBack_Enb),
	.sync_fast(sync_fast), .sync_jend(sync_jend), .SQSET(SQSET),
	.FAST_RST(FAST_RST), .TMODE(TMODE), .BypassDiv4(BypassDiv4),
	.tst_buferr(tst_buferr), .UTM_CHKERR(UTM_CHKERR),
	.FastStart(FastStart), .TEST_EYE_EN(TEST_EYE_EN),
	.FORCE_CRCERR(FORCE_CRCERR), .DIS_NARROW_SOF(DIS_NARROW_SOF),
	.RxDataOut_A(RxDataOut_A), .SquelchOut_A(SquelchOut_A),
	.DisconnectOut_A(DisconnectOut_A), .TERM_ON_A(TERM_ON_A),
	.RxDataOut_B(RxDataOut_B), .SquelchOut_B(SquelchOut_B),
        .DisconnectOut_B(DisconnectOut_B), .TERM_ON_B(TERM_ON_B),
	.RxDataOut_C(RxDataOut_C), .SquelchOut_C(SquelchOut_C),
        .DisconnectOut_C(DisconnectOut_C), .TERM_ON_C(TERM_ON_C),
	.RxDataOut_D(RxDataOut_D), .SquelchOut_D(SquelchOut_D),
        .DisconnectOut_D(DisconnectOut_D), .TERM_ON_D(TERM_ON_D),
	.RxDataOut_E(RxDataOut_E), .SquelchOut_E(SquelchOut_E),
        .DisconnectOut_E(DisconnectOut_E), .TERM_ON_E(TERM_ON_E),
	.RxDataOut_F(RxDataOut_F), .SquelchOut_F(SquelchOut_F),
        .DisconnectOut_F(DisconnectOut_F), .TERM_ON_F(TERM_ON_F),
	.RxDataOut_G(RxDataOut_G), .SquelchOut_G(SquelchOut_G),
        .DisconnectOut_G(DisconnectOut_G), .TERM_ON_G(TERM_ON_G),
	.RxDataOut_H(RxDataOut_H), .SquelchOut_H(SquelchOut_H),
        .DisconnectOut_H(DisconnectOut_H), .TERM_ON_H(TERM_ON_H),
	.DIS_TERM_ON_A(DIS_TERM_ON_A), .DIS_TERM_ON_B(DIS_TERM_ON_B),
	.DIS_TERM_ON_C(DIS_TERM_ON_C), .DIS_TERM_ON_D(DIS_TERM_ON_D),
	.DIS_TERM_ON_E(DIS_TERM_ON_E), .DIS_TERM_ON_F(DIS_TERM_ON_F),
	.DIS_TERM_ON_G(DIS_TERM_ON_G), .DIS_TERM_ON_H(DIS_TERM_ON_H),
	.autochk(autochk), .SetPowner_Dis(SetPowner_Dis),
	.PdPHY_Dis(PdPHY_Dis), .HsEnFB_Dis(HsEnFB_Dis),
	.USBLEGCTLSTS(USBLEGCTLSTS), .USBLEGSUP(USBLEGSUP),
	.PCI_R6AG(PCI_R6AG), .PCI_R6BG(PCI_R6BG), .PCI_R6CG(PCI_R6CG),
	.PCI_R6DG(PCI_R6DG), .PCI_R6FG(PCI_R6FG),
	.PCI_RBAR(PCI_RBAR), .PCI_RPCMD(PCI_RPCMD),
	//.PCI_R4EG(PCI_R4EG), .PCI_R4FG(PCI_R4FG),
	/*.EEMWR(EEMWR), .EEPRUN(EEPRUN), .EEPBUSY(EEPBUSY),
	.EEP_ADDR(EEP_ADDR), //.EEP_WDATA(EEP_WDATA),
	.EEP_RDATA(EEP_RDATA),*/ .SUBIDWE(SUBIDWE),
	.DISPDRCV(DISPDRCV), .CLKOFF_EN(CLKOFF_EN), .TXTMOUT_EN(TXTMOUT_EN),
	.TXDELAY_EN(TXDELAY_EN), .TXDELAY_PARM(TXDELAY_PARM),
	.TURN_PARM(TURN_PARM),
	.ENUSB1(ENUSB1), .ENUSB2(ENUSB2), .ENUSB3(ENUSB3), .ENUSB4(ENUSB4),
	.DIS_SOF_RUN(DIS_SOF_RUN), .SLEEPTIME_SEL(SLEEPTIME_SEL),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_WR(SRAM_WR), .SRAM_RUN(SRAM_RUN),
        .SRAM_RDATA1(SRAM_RDATA1), .SRAM_RDATA2(SRAM_RDATA2),
        .SRAM_RDATA3(SRAM_RDATA3), .SRAM_RDATA4(SRAM_RDATA4),
	.EN_DBG_PORT(EN_DBG_PORT) );
/*
    EEPCTL EEPCTL ( .EEPA7I(EEPA7I), .EEPA6I(EEPA6I), .EEPA5I(EEPA5I),
	.EEPA4I(EEPA4I), .EEPA3I(EEPA3I), .EEPA2I(EEPA2I),
	.EECBE(EECBE), .EEADO(EEADO), .EEPHASE(EEPHASE),
	.EIN15(EIN15), .EIN14(EIN14), .EIN13(EIN13), .EIN12(EIN12),
	.EIN11(EIN11), .EIN10(EIN10), .EIN9(EIN9), .EIN8(EIN8),
	.EIN7(EIN7), .EIN6(EIN6), .EIN5(EIN5), .EIN4(EIN4),
	.EIN3(EIN3), .EIN2(EIN2), .EIN1(EIN1), .EIN0(EIN0),
	.EEADDR5(EEADDR5), .EEADDR4(EEADDR4), .EEADDR3(EEADDR3),
	.EEADDR2(EEADDR2), .EEADDR1(EEADDR1), .EEADDR0(EEADDR0),
	.EEPBUSY(EEPBUSY), .EESTART(EESTART), .EECFGW0(EECFGW0),
	.EECFGW1(EECFGW1), .EECFGW2(EECFGW2),
	.EEPO15(EEPO15), .EEPO14(EEPO14), .EEPO13(EEPO13),
	.EEPO12(EEPO12), .EEPO11(EEPO11), .EEPO10(EEPO10),
	.EEPO9(EEPO9), .EEPO8(EEPO8), .EEPO7(EEPO7), .EEPO6(EEPO6),
	.EEPO5(EEPO5), .EEPO4(EEPO4), .EEPO3(EEPO3), .EEPO2(EEPO2),
	.EEPO1(EEPO1), .EEPO0(EEPO0), .EEPRUN(EEPRUN), .EEP_ADDR(EEP_ADDR),
	.LADO(LADO), .EEP_RDATA(EEP_RDATA),
	.PCI_R4EG(PCI_R4EG), .PCI_R4FG(PCI_R4FG),
	.WCOMPL(WCOMPL), .RCOMPL(RCOMPL), .PCICLK(PCICLK), .HRST_(HRST_) );

    EEPACCESS EEPACCESS ( .CS(EECS), .SK(EESK), .DI(EEDI), .EEDOG(EEDO),
	.EEPO15(EEPO15), .EEPO14(EEPO14), .EEPO13(EEPO13),
        .EEPO12(EEPO12), .EEPO11(EEPO11), .EEPO10(EEPO10),
        .EEPO9(EEPO9), .EEPO8(EEPO8), .EEPO7(EEPO7), .EEPO6(EEPO6),
        .EEPO5(EEPO5), .EEPO4(EEPO4), .EEPO3(EEPO3), .EEPO2(EEPO2),
        .EEPO1(EEPO1), .EEPO0(EEPO0), .WCOMPL(WCOMPL), .RCOMPL(RCOMPL),
	.EIN15(EIN15), .EIN14(EIN14), .EIN13(EIN13), .EIN12(EIN12),
	.EIN11(EIN11), .EIN10(EIN10), .EIN9(EIN9), .EIN8(EIN8),
	.EIN7(EIN7), .EIN6(EIN6), .EIN5(EIN5), .EIN4(EIN4),
	.EIN3(EIN3), .EIN2(EIN2), .EIN1(EIN1), .EIN0(EIN0), .EEADDR6(1'b0),
	.EEADDR5(EEADDR5), .EEADDR4(EEADDR4), .EEADDR3(EEADDR3),
	.EEADDR2(EEADDR2), .EEADDR1(EEADDR1), .EEADDR0(EEADDR0),
	.CISREAD(1'b0), .RDOPT(1'b0), .OHCIREAD(1'b0), .DPM(1'b0),
	.EEOPT(1'b0), .EEMWR(EEMWR), .EESTART(EESTART),
	.SYSCLK(PCICLK), .HRSTEZ(HRST_) );

    EEPMUX EEPMUX ( .ULADO(ULADO), .EEADO(EEADO), .LADO(LADO),
	.ULCBE(ULCBE), .EECBE(EECBE), .LCBE(LCBE),
	.UCFGW(UCFGW), .EECFGW(EECFGW2), .CFGW(CFGW), .EEPHASE(EEPHASE),
	.UPA7I(UPA7I), .UPA6I(UPA6I), .UPA5I(UPA5I), .UPA4I(UPA4I),
	.UPA3I(UPA3I), .UPA2I(UPA2I), .EEPA7I(EEPA7I), .EEPA6I(EEPA6I),
	.EEPA5I(EEPA5I), .EEPA4I(EEPA4I), .EEPA3I(EEPA3I),
	.EEPA2I(EEPA2I), .PA7I(PA7I), .PA6I(PA6I), .PA5I(PA5I),
	.PA4I(PA4I), .PA3I(PA3I), .PA2I(PA2I) );
*/
//wire [1:0] FRLSTSIZE;
//wire [31:0] ASYNCLISTADDR;

    HS_OPREG HS_OPREG ( .REGD31(REGD31), .REGD30(REGD30), .REGD29(REGD29), 
	.REGD28(REGD28), .REGD27(REGD27), .REGD26(REGD26), .REGD25(REGD25), 
	.REGD24(REGD24), .REGD23(REGD23), .REGD22(REGD22), .REGD21(REGD21), 
	.REGD20(REGD20), .REGD19(REGD19), .REGD18(REGD18), .REGD17(REGD17), 
	.REGD16(REGD16), .REGD15(REGD15), .REGD14(REGD14), .REGD13(REGD13), 
	.REGD12(REGD12), .REGD11(REGD11), .REGD10(REGD10), .REGD9(REGD9), 
	.REGD8(REGD8), .REGD7(REGD7), .REGD6(REGD6), .REGD5(REGD5), .REGD4(
	REGD4), .REGD3(REGD3), .REGD2(REGD2), .REGD1(REGD1), .REGD0(REGD0), 
	.ConfigFlag(ConfigFlag), .LIGHTRST(LIGHTRST), .ASYNC_EN(ASYNC_EN),
	.PERIOD_EN(PERIOD_EN), .FRLSTSIZE(FRLSTSIZE),
	.HCRESET(HCRESET), .RUN(RUN), .FLBASE(FLBASE), .RUN_C(RUN_C),
	.WR_FRNUM(WR_FRNUM), .ASYNCLISTADDR(ASYNCLISTADDR),
	.WR_ASYNCADDR(WR_ASYNCADDR), .FRNUM(FRNUM), .MAC_EOT(MAC_EOT),
	.MABORTS(MABORTS), .TABORTR(TABORTR), .RECLAMATION(RECLAMATION),
	.ASYNC_ACT(ASYNC_ACT), .PERIOD_ACT(PERIOD_ACT),
	.ROLLOVER_S(ROLLOVER_S), .UINTOE_(UINTOE_),
	.PORTCHG_S(PORTCHG_S), .DBGIRQ(DBGIRQ), .UIRQACT(UIRQACT),
	.INTR_DIS(INTR_DIS),
	.AD31I(LADO[31]), .AD30I(LADO[30]), 
	.AD29I(LADO[29]), .AD28I(LADO[28]), .AD27I(LADO[27]), .AD26I(LADO[26]),
	.AD25I(LADO[25]), .AD24I(LADO[24]), .AD23I(LADO[23]), .AD22I(LADO[22]),
	.AD21I(LADO[21]), .AD20I(LADO[20]), .AD19I(LADO[19]), 
	.AD18I(LADO[18]), .AD17I(LADO[17]), .AD16I(LADO[16]), .AD15I(LADO[15]),
	.AD14I(LADO[14]), .AD13I(LADO[13]), .AD12I(LADO[12]), .AD11I(
	LADO[11]), .AD10I(LADO[10]), .AD9I(LADO[9]), .AD8I(LADO[8]), .AD7I(
	LADO[7]), .AD6I(LADO[6]), .AD5I(LADO[5]), .AD4I(LADO[4]), .AD3I(
	LADO[3]), .AD2I(LADO[2]), .AD1I(LADO[1]), .AD0I(LADO[0]), /*.FRNUM15(
	FRNUM[15]), .FRNUM14(FRNUM[14]), .FRNUM13(FRNUM[13]), .FRNUM12(
	FRNUM[12]), .FRNUM11(FRNUM[11]), .FRNUM10(FRNUM[10]), .FRNUM9(FRNUM[9]
	), .FRNUM8(FRNUM[8]), .FRNUM7(FRNUM[7]), .FRNUM6(FRNUM[6]), .FRNUM5(
	FRNUM[5]), .FRNUM4(FRNUM[4]), .FRNUM3(FRNUM[3]), .FRNUM2(FRNUM[2]), 
	.FRNUM1(FRNUM[1]), .FRNUM0(FRNUM[0]), .HCHALT_S(HCHALT_S),*/
	.EHCI_IDLE(EHCI_IDLE), .HCHALT(HCHALT), .HSERR_S(HSERR_S),
	.ERRINT_S(ERRINT_S), .USBINT_S(USBINT_S), .USBINT(USBINT),
 	/*.HCERR_EN(HCERR),*/ .ERRINT_EN(ERRINT_EN), .USBINT_EN(USBINT_EN),
	.INTTHRESHOLD(INTTHRESHOLD), /*.IOCSPDINT(IOCSPDINT),
	.USBERRINT(USBERRINT),*/ .ERRINT(ERRINT), .INTASYNC_EN(INTASYNC_EN),
	.INTDOORBELL(INTDOORBELL), .INTASYNC_S(INTASYNC_S),
	.ASYNCINT(ASYNCINT), .INTASYNC(INTASYNC), .CMDRST_(CMDRST_),
	.PWR_STATE_D0(PWR_STATE_D0),

	/*.CONN1(CONN1), .CONN2(CONN2), .CONNCHG1(CONNCHG1), 
	.SDP1(SDP1), .SDP2(SDP2), .SDN1(SDN1), .SDN2(SDN2), */
	.PORTSC1(PORTSC1), .PORTSC2(PORTSC2), .PORTSC3(PORTSC3),
	.PORTSC4(PORTSC4), .PORTSC5(PORTSC5), .PORTSC6(PORTSC6),
	.PORTSC7(PORTSC7), .PORTSC8(PORTSC8),
	.CFG_CS(CFG_CS),
	.PSC_CBE2_A(PSC_CBE2_A), .PSC_CBE1_A(PSC_CBE1_A),
	.PSC_CBE0_A(PSC_CBE0_A),
 	.PSC_CBE2_B(PSC_CBE2_B), .PSC_CBE1_B(PSC_CBE1_B),
 	.PSC_CBE0_B(PSC_CBE0_B),
 	.PSC_CBE2_C(PSC_CBE2_C), .PSC_CBE1_C(PSC_CBE1_C),
 	.PSC_CBE0_C(PSC_CBE0_C),
 	.PSC_CBE2_D(PSC_CBE2_D), .PSC_CBE1_D(PSC_CBE1_D),
 	.PSC_CBE0_D(PSC_CBE0_D),
 	.PSC_CBE2_E(PSC_CBE2_E), .PSC_CBE1_E(PSC_CBE1_E),
 	.PSC_CBE0_E(PSC_CBE0_E),
 	.PSC_CBE2_F(PSC_CBE2_F), .PSC_CBE1_F(PSC_CBE1_F),
 	.PSC_CBE0_F(PSC_CBE0_F),
 	.PSC_CBE2_G(PSC_CBE2_G), .PSC_CBE1_G(PSC_CBE1_G),
 	.PSC_CBE0_G(PSC_CBE0_G),
 	.PSC_CBE2_H(PSC_CBE2_H), .PSC_CBE1_H(PSC_CBE1_H),
 	.PSC_CBE0_H(PSC_CBE0_H),
	.CBE3I_(LCBE[3]), .CBE2I_(LCBE[2]), 
	.CBE1I_(LCBE[1]), .CBE0I_(LCBE[0]), .REGW(REGW), .PA7I(PA7I), .PA6I(
	PA6I), .PA5I(PA5I), .PA4I(PA4I), .PA3I(PA3I), .PA2I(PA2I), 
	/*.OC1I_(OC1I_), .OC2I_(OC2I_),*/
	.PCICLK(PCICLK), .PCICLK_FREE(PCICLK_FREE), .HRST_(HRST_),
	.TEST_FORCE_ENABLE(TEST_FORCE_ENABLE), .ATPG_ENI(ATPG_ENI),
	.USBLEGCTLSTS(USBLEGCTLSTS), .USBLEGSUP(USBLEGSUP),
	.PCI_R6AG(PCI_R6AG), .PCI_R6BG(PCI_R6BG), .PCI_R6CG(PCI_R6CG),
	.PCI_R6DG(PCI_R6DG), .PCI_R6FG(PCI_R6FG),
	.PCI_RBAR(PCI_RBAR), .PCI_RPCMD(PCI_RPCMD), .USMIO(USMIO),
	.SUBIDWE(SUBIDWE),
	.ENUSB1(ENUSB1), .ENUSB2(ENUSB2), .ENUSB3(ENUSB3), .ENUSB4(ENUSB4),
	.DIS_SOF_RUN(DIS_SOF_RUN), .UTM_RUN(UTM_RUN),
	.FRNUM_PCLK_LATCH_66(FRNUM_PCLK_LATCH_66),
	.EN_DBG_PORT(EN_DBG_PORT),
	.DBGPORT_R00G(DBGPORT_R00G), .DBGPORT_R01G(DBGPORT_R01G),
	.DBGPORT_R02G(DBGPORT_R02G), .DBGPORT_R03G(DBGPORT_R03G),
        .DBGPORT_R04G(DBGPORT_R04G), .DBGPORT_R05G(DBGPORT_R05G),
	.DBGPORT_R08G(DBGPORT_R08G), .DBGPORT_R09G(DBGPORT_R09G),
        .DBGPORT_R0AG(DBGPORT_R0AG), .DBGPORT_R0BG(DBGPORT_R0BG),
	.DBGPORT_R0CG(DBGPORT_R0CG), .DBGPORT_R0DG(DBGPORT_R0DG),
        .DBGPORT_R0EG(DBGPORT_R0EG), .DBGPORT_R0FG(DBGPORT_R0FG),
	.DBGPORT_R10G(DBGPORT_R10G), .DBGPORT_R11G(DBGPORT_R11G),
        .DBGPORT_SC(DBGPORT_SC), .DBGPORT_PID(DBGPORT_PID),
	.DBGPORT_ADDR(DBGPORT_ADDR),
        .DBGPORT_BUF1(DBGPORT_BUF1), .DBGPORT_BUF2(DBGPORT_BUF2) );

    HS_DBG_OPREG HS_DBG_OPREG ( .ADI(LADO), .EN_DBG_PORT(EN_DBG_PORT),
	.DBGPORT_R00G(DBGPORT_R00G), .DBGPORT_R01G(DBGPORT_R01G),
        .DBGPORT_R02G(DBGPORT_R02G), .DBGPORT_R03G(DBGPORT_R03G),
        .DBGPORT_R04G(DBGPORT_R04G), .DBGPORT_R05G(DBGPORT_R05G),
        .DBGPORT_R10G(DBGPORT_R10G), .DBGPORT_R11G(DBGPORT_R11G),
        .DBGPORT_SC(DBGPORT_SC), .DBGPORT_PID(DBGPORT_PID),
	.DBGPORT_ADDR(DBGPORT_ADDR),
        .DBG_COMPL(DBG_COMPL), .DBG_XACTERR(DBG_XACTERR),
	.PORT_SUSPEND(PORTSC1[7]), .PORT_RESET(PORTSC1[8]),
        .DBG_RXBCNT(DBG_RXBCNT), .DBG_RXPID(DBG_RXPID),
	.DBG_ENABLE_WC(DBG_ENABLE_WC), .PORT_ENDIS(PORTSC1[2]),
        .PCICLK(PCICLK), .PCICLK_FREE(PCICLK_FREE), .CMDRST_(CMDRST_) );

    UTGTCTL UTGTCTL ( .THIT(THIT), .ADRG(ADRG), .ADS(UADS), .TADOE(TADOE), .TERM(
	TERM), /*.RDYACK(RDYACK),*/ .FRAME0(FRAME0), .FRAME4(FRAME4), .TDATA(TDATA
	), .TRDYO_(TRDYO_), .STOPO_(STOPO_), .DEVSELO_(DEVSELO_), .TRDYOE_(
	TRDYOE_), .TPAROE_(TPAROE_), .IRDYI_(IRDYI_), .DEVSELI_(DEVSELI_), 
	.FRAMEI_(FRAMEI_), .TRDYI_(TRDYI_), .DEVS0(DEVS0), .HIT(UHIT), .LRDY(
	ULRDY), .TGWR(LCMD0), .HITKBC(1'b0),
	.PCICLK(PCICLK_FREE), .HRST_(HRST_), .PCIS_ACT(PCIS_ACT),
	.ADS_PRE(ADS_PRE), .PMSTR(PMSTR), .TRDYOED_(TRDYOED_),
	.ATPG_EN(ATPG_ENI) );
    ziva rev7 ( .A(GND), .Y(REVID7) );
    ziva rev6 ( .A(VDD), .Y(REVID6) );
    ziva rev5 ( .A(VDD), .Y(REVID5) );
    ziva rev4 ( .A(GND), .Y(REVID4) );
    ziva rev3 ( .A(VDD), .Y(REVID3) );
    ziva rev2 ( .A(VDD), .Y(REVID2) );
    ziva rev1 ( .A(VDD), .Y(REVID1) );
    ziva rev0 ( .A(VDD), .Y(REVID0) );
    /*ziva usb7 ( .A(VDD), .Y(USBSPEC7) );
    ziva usb6 ( .A(VDD), .Y(USBSPEC6) );
    ziva usb5 ( .A(GND), .Y(USBSPEC5) );
    ziva usb4 ( .A(VDD), .Y(USBSPEC4) );
    ziva usb3 ( .A(VDD), .Y(USBSPEC3) );
    ziva usb2 ( .A(VDD), .Y(USBSPEC2) );
    ziva usb1 ( .A(VDD), .Y(USBSPEC1) );
    ziva usb0 ( .A(VDD), .Y(USBSPEC0) );*/
    ziva mlat7 ( .A(VDD), .Y(MAXLAT7) );
    ziva mlat6 ( .A(VDD), .Y(MAXLAT6) );
    ziva mlat5 ( .A(VDD), .Y(MAXLAT5) );
    ziva mlat4 ( .A(VDD), .Y(MAXLAT4) );
    ziva mlat3 ( .A(VDD), .Y(MAXLAT3) );
    ziva mlat2 ( .A(VDD), .Y(MAXLAT2) );
    ziva mlat1 ( .A(VDD), .Y(MAXLAT1) );
    ziva mlat0 ( .A(VDD), .Y(MAXLAT0) );
    ziva mgnt7 ( .A(VDD), .Y(MINGNT7) );
    ziva mgnt6 ( .A(VDD), .Y(MINGNT6) );
    ziva mgnt5 ( .A(VDD), .Y(MINGNT5) );
    ziva mgnt4 ( .A(VDD), .Y(MINGNT4) );
    ziva mgnt3 ( .A(VDD), .Y(MINGNT3) );
    ziva mgnt2 ( .A(VDD), .Y(MINGNT2) );
    ziva mgnt1 ( .A(VDD), .Y(MINGNT1) );
    ziva mgnt0 ( .A(VDD), .Y(MINGNT0) );
endmodule


module HS_FFCTL ( USBDAT, HOSTDAT, LATCHDAT, USBPOP, CLK60M, BUISTRT, WPR0, 
    WPR1, EOT, PCICLK, ADI, FPUSH, FPOP, MDO, MDI, WMA, RMA, PCIWRT, PCIREAD, 
    RXFIFO, UCBEO_, RXSTRT, XMITSTRT, FIFO_OK, FFRDPCI, FBE_, TDMAEND, RDMAEND, 
    RXPKTEND, TRST_, FCOUNT, FFULL, FEMPTY, RXERR, TEST_PACKET, TESTAD, 
    TESTDOUT, TESTPKTOK, ATPG_ENI );
input  [7:0] USBDAT;
output [7:0] HOSTDAT;
input  [31:0] ADI;
input  [31:0] MDO;
output [8:0] WMA;
input  [3:0] UCBEO_;
output [8:0] FCOUNT;
output [3:0] FBE_;
output [31:0] FFRDPCI;
output [31:0] MDI;
output [8:0] RMA;
output [3:0] TESTAD;
input  [31:0] TESTDOUT;
input  LATCHDAT, USBPOP, CLK60M, BUISTRT, WPR0, WPR1, EOT, PCICLK, PCIWRT, 
    PCIREAD, RXFIFO, RXSTRT, XMITSTRT, TDMAEND, RDMAEND, TRST_, RXERR, 
    TEST_PACKET, ATPG_ENI;
output FPUSH, FPOP, FIFO_OK, RXPKTEND, FFULL, FEMPTY, TESTPKTOK;
    wire USBFFTMP_12, N_FIFOCNT_8, FPOP_T1737, PCIWRT_TEST, FIFOCNT_2, 
        FFRDUSB2141_7, FFRDUSB_13, PCIDATA_T1208_11, FFRDUSB2141_13, 
        FFRDPCI1761_9, USBFFTMP655_16, SPAREO6, USBFFTMP655_31, c1328_7, 
        PCIDATA_T1208_9, USBFFTMP_9, FFRDPCI1761_22, FSIZE1570_0, PIPE_START_T, 
        PCIDATA_23, PCIDATA_T_21, PSH, PCIDATA_7, rptr_7, END_BE_1, 
        USBTMP396_6, FFRDUSB_4, USBTMP396_22, N_FIFOCNT_1, USBTMP396_17, 
        EOT3_T, USBTMP396_30, n_rptr_7, PCIDATA_T_14, PCIDATA_T1208_18, 
        USBFFTMP655_5, PCIDATA_16, PCIDATA_31, wptr_4, EOT3_T1447, 
        FFRDPCI1761_17, FFRDPCI1761_30, FFRDPCI1761_0, PCIDATA_T_7, 
        PCIDATA_T1208_0, USBFFTMP655_23, N_FIFOCNT835_6, PCIDATA_T_28, 
        PCIDATA_T1208_24, FFRDUSB_26, FFRDUSB2141_26, USBFFTMP_0, USBFFTMP_27, 
        END_BE2076_1, TESTAD1135_1, PCIDATA_9, USBTMP396_8, USBFFTMP_20, 
        c1328_9, USBFFTMP655_24, N_FIFOCNT835_1, PCIDATA_T1208_7, PCIDATA_T_0, 
        USBFFTMP_7, SPAREO0_, FFRDUSB2141_21, FFRDUSB_21, PCIDATA_T1208_23, 
        FFRDUSB2141_9, USBFFTMP655_2, PCIDATA_11, PCIDATA_T_13, FFRDPCI1761_7, 
        USBFFTMP655_18, SPAREO8, wptr_3, FFRDPCI1761_10, n_rptr_0, 
        USBTMP396_10, N_FIFOCNT_6, EOT_PCLK_T, TESTAD1143_1, FFRDUSB_3, 
        USBTMP396_1, rptr_0, PCIDATA_0, FBE_2296_1, USBTMP396_25, USBFFTMP_29, 
        FFRDPCI1761_25, PCIDATA_T_9, N_FIFOCNT835_8, PCIDATA_T_26, FFRDUSB_28, 
        FFRDUSB2141_28, PCIDATA_24, PIPE_START1493, TCNT1958_0, FFRDUSB2141_14, 
        PCIDATA_T1208_16, FFRDUSB_14, PCIDATA_18, FFRDUSB2141_0, 
        PCIDATA_T1208_31, FFRDPCI1761_19, USBFFTMP655_11, SPAREO1, FSIZE_1, 
        USBTMP396_19, USBFFTMP_15, TEST_START, RDFF_EQ_WAIT, FIFOCNT_5, 
        n_rptr_1, USBTMP396_11, N_FIFOCNT_7, FPUSH770, FFRDUSB2141_8, 
        PCIDATA_10, USBFFTMP655_3, PCIDATA_T_12, FFRDPCI1761_6, USBFFTMP655_19, 
        SPAREO9, wptr_2, EOT3_2T, FFRDPCI1761_11, c1328_8, PCIDATA_T1208_6, 
        USBFFTMP655_25, N_FIFOCNT835_0, PCIDATA_T_1, LDWPR, USBFFTMP_6, 
        FFRDUSB_20, PCIDATA_T1208_22, FFRDUSB2141_20, rptr_8, PCIDATA_8, 
        USBTMP396_9, USBFFTMP_21, PROCESS, LDWPR2000, USBTMP396_18, FSIZE_0, 
        USBFFTMP_14, n_rptr_8, EOT_T, FIFOCNT_4, val628_1, PCIWRT_TEST1184, 
        PCIDATA_T1208_17, FFRDUSB_15, TCNT1958_1, FFRDUSB2141_15, PCIDATA_19, 
        FFRDUSB2141_1, PCIDATA_T1208_30, FFRDPCI1761_18, FIFO_OK1699, 
        USBFFTMP655_10, SPAREO0, EOT_2T, FFRDPCI1761_24, PCIDATA_T_8, 
        PROCESS2334, FPOP_ONCE, c1328_1, FFRDUSB2141_29, FFRDUSB_29, 
        PCIDATA_T_27, PCIDATA_25, FFRDUSB_2, TESTAD1143_0, USBTMP396_0, 
        PCIDATA_1, rptr_1, FBE_2296_0, USBTMP396_24, USBFFTMP_28, rptr_6, 
        PCIDATA_6, USBTMP396_7, END_BE_0, FFRDUSB_5, USBTMP396_23, c1328_6, 
        PCIDATA_T1208_8, FFRDPCI1761_23, FSIZE1570_1, USBFFTMP_8, PCIDATA_22, 
        PCIDATA_T_20, FFRDUSB2141_6, RXPKTEND2408, FFRDUSB2141_12, FFRDUSB_12, 
        PCIDATA_T1208_10, FFRDPCI1761_8, SPAREO7, USBFFTMP655_17, 
        USBFFTMP655_30, FPOP_ONCE1612, USBFFTMP_13, PIPE_START_2T, FIFOCNT_3, 
        USBFFTMP_26, END_BE2076_0, PCIDATA_T_6, USBFFTMP655_22, N_FIFOCNT835_7, 
        PCIDATA_T1208_1, FFRDUSB2141_27, PCIDATA_T1208_25, PCIDATA_T_29, 
        FFRDUSB_27, USBFFTMP_1, PCIDATA_T_15, PCIDATA_T1208_19, PCIDATA_17, 
        USBFFTMP655_4, PCIDATA_30, FFRDPCI1761_16, wptr_5, FFRDPCI1761_31, 
        FFRDPCI1761_1, N_FIFOCNT_0, USBTMP396_16, USBTMP396_31, n_rptr_6, 
        RDFFNXT_1, FIFOCNT_1, PSH1244, USBFFTMP_11, SPAREO5, USBFFTMP655_15, 
        FFRDUSB_10, PCIDATA_T1208_12, FFRDUSB2141_10, FFRDUSB2141_4, 
        PCIDATA_20, PCIDATA_T_22, FFRDPCI1761_21, USBFFTMP655_29, c1328_4, 
        USBTMP396_21, ST_BE_0, ST_BE2037_1, END_BE_2, USBTMP396_5, FFRDUSB_7, 
        rptr_4, PCIDATA_4, FIFOCNT_8, RCNT351_1, USBFFTMP_18, FSIZE1554_1, 
        n_rptr_4, N_FIFOCNT_2, USBTMP396_14, wptr_7, FFRDPCI1761_3, 
        FFRDPCI1761_14, PCIDATA_T_30, FFRDUSB2141_19, PCIDATA_T_17, FFRDUSB_19, 
        EOT_PCLK_2T, PCIDATA_15, USBFFTMP655_6, LDWPR_2T, RCNT_1, USBFFTMP_3, 
        FFRDUSB_25, PCIDATA_T1208_27, FFRDUSB2141_25, PCIDATA_29, 
        PCIDATA_T1208_3, USBFFTMP655_20, N_FIFOCNT835_5, FFRDPCI1761_28, 
        PCIDATA_T_4, END_BE2076_2, USBFFTMP_24, TESTAD1135_2, USBTMP396_28, 
        USBFFTMP_23, FFRDUSB_9, FFRDUSB2141_22, USBFFTMP_4, PCIDATA_T1208_20, 
        FFRDUSB_22, PCIDATA_T_3, USBFFTMP655_27, N_FIFOCNT835_2, 
        PCIDATA_T1208_4, FFRDPCI1761_13, wptr_0, FFRDPCI1761_4, PCIDATA_12, 
        USBFFTMP655_1, PCIDATA_T_10, RXWRT, USBTMP396_13, N_FIFOCNT_5, 
        n_rptr_3, USBTMP396_26, FIRSTDW2259, PCIDATA_3, rptr_3, FBE_2296_2, 
        FFRDUSB_0, TESTAD1143_2, USBTMP396_2, PCIDATA_T1208_29, PCIDATA_T_25, 
        PCIDATA_27, c1328_3, RCNT_0, FFRDPCI1761_26, USBFFTMP655_12, SPAREO2, 
        FFRDUSB2141_3, FFRDUSB_30, FFRDUSB2141_30, FFRDUSB2141_17, 
        PCIDATA_T_19, FFRDUSB_17, PCIDATA_T1208_15, USBFFTMP655_8, FIFOCNT_6, 
        UPOP, USBFFTMP_16, USBFFTMP_31, N_FIFOCNT_4, USBTMP396_12, n_rptr_2, 
        wptr_1, FFRDPCI1761_12, FFRDPCI1761_5, PCIDATA_13, USBFFTMP655_0, 
        PCIDATA_T_11, PCIDATA_T1208_21, FFRDUSB_23, LDWPR_T, FFRDUSB2141_23, 
        USBFFTMP_5, PCIDATA_T_2, PCIDATA_T1208_5, N_FIFOCNT835_3, 
        USBFFTMP655_26, USBFFTMP_22, FFRDUSB_8, USBREAD, FIFOCNT_7, 
        USBFFTMP_17, USBFFTMP_30, USBFFTMP655_13, SPAREO3, wptr_8, SPAREO1_, 
        FFRDUSB2141_2, FFRDUSB_31, PCIDATA_T_18, FPOP_T, FFRDUSB2141_31, 
        FFRDUSB_16, PCIDATA_T1208_14, FFRDUSB2141_16, USBFFTMP655_9, 
        PCIDATA_T1208_28, PCIDATA_T_24, PCIDATA_26, c1328_2, FFRDPCI1761_27, 
        USBTMP396_27, rptr_2, PCIDATA_2, FBE_2296_3, FFRDUSB_1, TESTAD1143_3, 
        USBTMP396_3, USBTMP396_20, USBTMP396_4, END_BE_3, ST_BE2037_0, 
        FFRDUSB_6, FIRSTDW, PCIDATA_5, rptr_5, RXPKTEND_T2371, PCIDATA_21, 
        PCIDATA_T_23, FFRDPCI1761_20, c1328_5, USBFFTMP655_28, USBFFTMP655_14, 
        SPAREO4, FFRDUSB2141_11, FFRDUSB_11, PCIDATA_T1208_13, FFRDUSB2141_5, 
        TCNT1929_1, RDFFNXT_0, FIFOCNT_0, RCNT322_1, USBFFTMP_10, TESTAD1135_3, 
        END_BE2076_3, USBFFTMP_25, USBTMP396_29, USBFFTMP_2, FFRDUSB2141_24, 
        FFRDUSB_24, PCIDATA_T1208_26, PCIDATA_28, N_FIFOCNT835_4, 
        USBFFTMP655_21, PCIDATA_T1208_2, FFRDPCI1761_29, PCIDATA_T_5, 
        PIPE_START, FFRDPCI1761_2, wptr_6, FFRDPCI1761_15, PCIDATA_T_31, 
        FFRDUSB_18, EOT_PCLK, PCIDATA_T_16, FFRDUSB2141_18, PCIDATA_14, 
        USBFFTMP655_7, RCNT351_0, USBFFTMP_19, n_rptr_5, FSIZE1554_0, 
        N_FIFOCNT_3, USBTMP396_15, n2586, n2587, n2949, n2951, n2952, n2953, 
        n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
        n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
        n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
        n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
        n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3003, n3004, 
        n3005, n3006, n3007, n3009, n3010, n3011, n3012, n3013, n3014, n3015, 
        n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, 
        n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, 
        n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, 
        n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, 
        n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
        add_416_carry_8, add_416_carry_6, add_416_carry_7, add_416_carry_2, 
        add_416_carry_5, add_416_carry_4, add_416_carry_3, add_536_carry_8, 
        add_536_carry_1, add_536_carry_7, add_536_carry_6, add_536_carry_2, 
        add_536_carry_5, add_536_carry_4, add_536_carry_3, add_362_carry_2, 
        add_362_carry_3, r255_carry_1, r235_carry_8, r235_carry_1, 
        r235_carry_7, r235_carry_6, r235_carry_2, r235_carry_5, r235_carry_4, 
        r235_carry_3, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, 
        n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, 
        n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, 
        n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, 
        n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, 
        n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, 
        n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, 
        n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, 
        n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, 
        n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, 
        n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, 
        n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, 
        n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, 
        n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, 
        n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, 
        n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, 
        n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, 
        n3232, n3233, _cell_531_U41_Z_0, _cell_531_U22_Z_0, n3234, n3235, 
        n3236, n3237;
    zivb SPARE697 ( .A(SPAREO4), .Y(SPAREO5) );
    zdffrb SPARE690 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE699 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE691 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE698 ( .A(SPAREO5), .Y(SPAREO6) );
    znr3b SPARE696 ( .A(SPAREO2), .B(n2961), .C(SPAREO0_), .Y(SPAREO4) );
    zoai21b SPARE694 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE693 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zaoi211b SPARE692 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE695 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zor2b U1102 ( .A(FIRSTDW2259), .B(n3191), .Y(n3219) );
    zxo2b U1103 ( .A(RCNT_0), .B(RCNT_1), .Y(RCNT322_1) );
    zor2b U1104 ( .A(RCNT_0), .B(n3101), .Y(n3134) );
    zor2b U1105 ( .A(n3075), .B(n3107), .Y(n3106) );
    zan2b U1106 ( .A(FPOP), .B(FPUSH), .Y(n3065) );
    zor2b U1107 ( .A(n3066), .B(n3105), .Y(n3198) );
    zivb U1108 ( .A(n3198), .Y(n3195) );
    zxo2b U1109 ( .A(n2586), .B(n2587), .Y(TCNT1929_1) );
    zmux21lb U1110 ( .A(n3218), .B(FSIZE_1), .S(FSIZE_0), .Y(n3203) );
    zao21b U1111 ( .A(EOT3_2T), .B(n3205), .C(PIPE_START), .Y(n3222) );
    zivb U1112 ( .A(n3097), .Y(n3095) );
    zmux21lb U1113 ( .A(n3191), .B(n3209), .S(n2998), .Y(TCNT1958_0) );
    zmux21lb U1114 ( .A(n2586), .B(n3190), .S(UPOP), .Y(n3209) );
    zmux21hb U1115 ( .A(TESTAD[0]), .B(n3183), .S(n2953), .Y(TESTAD1143_0) );
    zmux21lb U1116 ( .A(n3211), .B(n3214), .S(n2999), .Y(RCNT351_0) );
    zao22b U1117 ( .A(FIFOCNT_0), .B(n3088), .C(N_FIFOCNT835_0), .D(n2955), 
        .Y(N_FIFOCNT_0) );
    zmux21lb U1118 ( .A(n3146), .B(n2993), .S(n3006), .Y(USBTMP396_12) );
    zmux21lb U1119 ( .A(n3123), .B(n2972), .S(LATCHDAT), .Y(USBTMP396_30) );
    zmux21lb U1120 ( .A(n3142), .B(n2989), .S(n3006), .Y(USBTMP396_16) );
    zor2b U1121 ( .A(PCIREAD), .B(FIRSTDW), .Y(FIRSTDW2259) );
    zor2b U1122 ( .A(n3113), .B(n3077), .Y(n3078) );
    zivb U1123 ( .A(n3134), .Y(n3113) );
    zmux21lb U1124 ( .A(n2967), .B(n3154), .S(n3207), .Y(USBFFTMP655_6) );
    zmux21lb U1125 ( .A(n2978), .B(n3164), .S(n3207), .Y(USBFFTMP655_25) );
    zor2b U1126 ( .A(RCNT_0), .B(RCNT_1), .Y(n3079) );
    zivb U1127 ( .A(n3079), .Y(n3107) );
    zmux21lb U1128 ( .A(n2990), .B(n3175), .S(n3233), .Y(USBFFTMP655_15) );
    zmux21lb U1129 ( .A(n2977), .B(n3163), .S(n3233), .Y(USBFFTMP655_26) );
    zao21b U1130 ( .A(RXWRT), .B(_cell_531_U22_Z_0), .C(PSH), .Y(FPUSH770) );
    zmux21lb U1131 ( .A(n3204), .B(n3219), .S(n3202), .Y(n3069) );
    zao22b U1132 ( .A(END_BE_3), .B(n3071), .C(FBE_[3]), .D(n2959), .Y(
        FBE_2296_3) );
    zao22b U1133 ( .A(rptr_1), .B(n3084), .C(c1328_2), .D(n2956), .Y(n_rptr_1)
         );
    zhadrb add_416_U1_1_1 ( .A(rptr_1), .B(rptr_0), .CO(add_416_carry_2), .S(
        c1328_2) );
    zmux21lb U1134 ( .A(n3150), .B(n2997), .S(LATCHDAT), .Y(USBTMP396_0) );
    zmux21lb U1135 ( .A(n3108), .B(n2963), .S(LATCHDAT), .Y(USBTMP396_9) );
    zor2b U1136 ( .A(n2960), .B(FIFO_OK), .Y(FIFO_OK1699) );
    zmux21lb U1137 ( .A(n2986), .B(n3171), .S(n3233), .Y(USBFFTMP655_19) );
    zmux21lb U1138 ( .A(n2983), .B(n3168), .S(n3207), .Y(USBFFTMP655_21) );
    zmux21lb U1139 ( .A(n2991), .B(n3176), .S(n3207), .Y(USBFFTMP655_14) );
    zmux21lb U1140 ( .A(n2972), .B(n3158), .S(n3207), .Y(USBFFTMP655_30) );
    zmux21lb U1141 ( .A(n2995), .B(n3180), .S(n3207), .Y(USBFFTMP655_10) );
    zor2b U1142 ( .A(RXSTRT), .B(XMITSTRT), .Y(LDWPR2000) );
    zmux21lb U1143 ( .A(n3046), .B(n3034), .S(wptr_8), .Y(n3055) );
    zor2b U1144 ( .A(n3040), .B(n3017), .Y(n3046) );
    zmux21lb U1145 ( .A(n3040), .B(n3020), .S(wptr_7), .Y(n3056) );
    zmux21lb U1146 ( .A(n3047), .B(n3019), .S(wptr_6), .Y(n3057) );
    zor2b U1147 ( .A(n3039), .B(n3016), .Y(n3047) );
    zmux21lb U1148 ( .A(n3039), .B(n3048), .S(wptr_5), .Y(n3058) );
    zivb U1149 ( .A(n3045), .Y(n3048) );
    zao21b U1150 ( .A(n3099), .B(n3013), .C(n3044), .Y(n3045) );
    zmux21lb U1151 ( .A(n3049), .B(n3050), .S(wptr_4), .Y(n3059) );
    zor2b U1152 ( .A(n3038), .B(n3014), .Y(n3049) );
    zivb U1153 ( .A(n3044), .Y(n3050) );
    zao21b U1154 ( .A(n3099), .B(n3014), .C(n3043), .Y(n3044) );
    zmux21lb U1155 ( .A(n3038), .B(n3051), .S(wptr_3), .Y(n3060) );
    zivb U1156 ( .A(n3043), .Y(n3051) );
    zoai21b U1157 ( .A(wptr_2), .B(n3035), .C(n3018), .Y(n3043) );
    zmux21lb U1158 ( .A(n3052), .B(n3018), .S(wptr_2), .Y(n3061) );
    zor2b U1159 ( .A(n3037), .B(n3012), .Y(n3052) );
    zmux21lb U1160 ( .A(n3037), .B(n3053), .S(wptr_1), .Y(n3062) );
    zivb U1161 ( .A(n3041), .Y(n3053) );
    zoai21b U1162 ( .A(wptr_0), .B(n3035), .C(n3042), .Y(n3041) );
    zmux21lb U1163 ( .A(n3054), .B(n3042), .S(wptr_0), .Y(n3063) );
    zor2b U1164 ( .A(n3036), .B(n3035), .Y(n3054) );
    zivb U1165 ( .A(n3099), .Y(n3035) );
    zivb U1166 ( .A(n3036), .Y(n3042) );
    zor2b U1167 ( .A(FFULL), .B(_cell_531_U22_Z_0), .Y(n3036) );
    zmux21lb U1168 ( .A(n3210), .B(n3213), .S(n2999), .Y(RCNT351_1) );
    zmux21lb U1169 ( .A(n3122), .B(n2971), .S(LATCHDAT), .Y(USBTMP396_31) );
    zmux21lb U1170 ( .A(n3126), .B(n2974), .S(LATCHDAT), .Y(USBTMP396_29) );
    zmux21lb U1171 ( .A(n3136), .B(n2983), .S(n3006), .Y(USBTMP396_21) );
    zmux21lb U1172 ( .A(n3137), .B(n2984), .S(n3006), .Y(USBTMP396_20) );
    zmux21lb U1173 ( .A(n3139), .B(n2986), .S(n3006), .Y(USBTMP396_19) );
    zmux21lb U1174 ( .A(n3140), .B(n2987), .S(n3006), .Y(USBTMP396_18) );
    zmux21lb U1175 ( .A(n3141), .B(n2988), .S(n3006), .Y(USBTMP396_17) );
    zmux21lb U1176 ( .A(n3144), .B(n2991), .S(n3006), .Y(USBTMP396_14) );
    zmux21lb U1177 ( .A(n3148), .B(n2995), .S(n3006), .Y(USBTMP396_10) );
    zmux21lb U1178 ( .A(n3111), .B(n2964), .S(LATCHDAT), .Y(USBTMP396_8) );
    zmux21lb U1179 ( .A(n3116), .B(n2967), .S(LATCHDAT), .Y(USBTMP396_6) );
    zmux21lb U1180 ( .A(n3118), .B(n2968), .S(LATCHDAT), .Y(USBTMP396_5) );
    zmux21lb U1181 ( .A(n3120), .B(n2969), .S(LATCHDAT), .Y(USBTMP396_4) );
    zmux21lb U1182 ( .A(n3124), .B(n2973), .S(LATCHDAT), .Y(USBTMP396_3) );
    zmux21lb U1183 ( .A(n3138), .B(n2985), .S(n3006), .Y(USBTMP396_2) );
    zmux21lb U1184 ( .A(n2971), .B(n3157), .S(n3233), .Y(USBFFTMP655_31) );
    zmux21lb U1185 ( .A(n2974), .B(n3160), .S(n3207), .Y(USBFFTMP655_29) );
    zmux21lb U1186 ( .A(n2975), .B(n3161), .S(n3233), .Y(USBFFTMP655_28) );
    zmux21lb U1187 ( .A(n2976), .B(n3162), .S(n3207), .Y(USBFFTMP655_27) );
    zmux21lb U1188 ( .A(n2979), .B(n3165), .S(n3233), .Y(USBFFTMP655_24) );
    zmux21lb U1189 ( .A(n2981), .B(n3166), .S(n3207), .Y(USBFFTMP655_23) );
    zmux21lb U1190 ( .A(n2982), .B(n3167), .S(n3233), .Y(USBFFTMP655_22) );
    zivb U1191 ( .A(USBDAT[6]), .Y(n3117) );
    zmux21lb U1192 ( .A(n2984), .B(n3169), .S(n3233), .Y(USBFFTMP655_20) );
    zmux21lb U1193 ( .A(n2987), .B(n3172), .S(n3207), .Y(USBFFTMP655_18) );
    zmux21lb U1194 ( .A(n2988), .B(n3173), .S(n3233), .Y(USBFFTMP655_17) );
    zmux21lb U1195 ( .A(n2989), .B(n3174), .S(n3207), .Y(USBFFTMP655_16) );
    zmux21lb U1196 ( .A(n2992), .B(n3177), .S(n3233), .Y(USBFFTMP655_13) );
    zmux21lb U1197 ( .A(n2993), .B(n3178), .S(n3207), .Y(USBFFTMP655_12) );
    zmux21lb U1198 ( .A(n2994), .B(n3179), .S(n3233), .Y(USBFFTMP655_11) );
    zmux21lb U1199 ( .A(n2963), .B(n3151), .S(n3233), .Y(USBFFTMP655_9) );
    zmux21lb U1200 ( .A(n2964), .B(n3152), .S(n3207), .Y(USBFFTMP655_8) );
    zmux21lb U1201 ( .A(n2966), .B(n3153), .S(n3233), .Y(USBFFTMP655_7) );
    zivb U1202 ( .A(USBDAT[7]), .Y(n3115) );
    zmux21lb U1203 ( .A(n2968), .B(n3155), .S(n3233), .Y(USBFFTMP655_5) );
    zivb U1204 ( .A(USBDAT[5]), .Y(n3119) );
    zmux21lb U1205 ( .A(n2969), .B(n3156), .S(n3207), .Y(USBFFTMP655_4) );
    zivb U1206 ( .A(USBDAT[4]), .Y(n3121) );
    zmux21lb U1207 ( .A(n2973), .B(n3159), .S(n3233), .Y(USBFFTMP655_3) );
    zivb U1208 ( .A(USBDAT[3]), .Y(n3125) );
    zmux21lb U1209 ( .A(n2985), .B(n3170), .S(n3207), .Y(USBFFTMP655_2) );
    zivb U1210 ( .A(USBDAT[2]), .Y(n3130) );
    zmux21lb U1211 ( .A(n2996), .B(n3181), .S(n3233), .Y(USBFFTMP655_1) );
    zivb U1212 ( .A(USBDAT[1]), .Y(n3109) );
    zmux21lb U1213 ( .A(n2997), .B(n3182), .S(n3207), .Y(USBFFTMP655_0) );
    zivb U1214 ( .A(USBDAT[0]), .Y(n3112) );
    zao22b U1215 ( .A(FIFOCNT_8), .B(n3088), .C(N_FIFOCNT835_8), .D(n2955), 
        .Y(N_FIFOCNT_8) );
    zxo3b r235_U1_8 ( .A(FIFOCNT_8), .B(_cell_531_U22_Z_0), .C(r235_carry_8), 
        .Y(N_FIFOCNT835_8) );
    zao22b U1216 ( .A(FIFOCNT_7), .B(n3088), .C(N_FIFOCNT835_7), .D(n2955), 
        .Y(N_FIFOCNT_7) );
    zao22b U1217 ( .A(FIFOCNT_6), .B(n3088), .C(N_FIFOCNT835_6), .D(n2955), 
        .Y(N_FIFOCNT_6) );
    zao22b U1218 ( .A(FIFOCNT_5), .B(n3088), .C(N_FIFOCNT835_5), .D(n2955), 
        .Y(N_FIFOCNT_5) );
    zao22b U1219 ( .A(FIFOCNT_4), .B(n3088), .C(N_FIFOCNT835_4), .D(n2955), 
        .Y(N_FIFOCNT_4) );
    zao22b U1220 ( .A(FIFOCNT_3), .B(n3088), .C(N_FIFOCNT835_3), .D(n2955), 
        .Y(N_FIFOCNT_3) );
    zao22b U1221 ( .A(FIFOCNT_2), .B(n3088), .C(N_FIFOCNT835_2), .D(n2955), 
        .Y(N_FIFOCNT_2) );
    zao22b U1222 ( .A(FIFOCNT_1), .B(n3088), .C(N_FIFOCNT835_1), .D(n2955), 
        .Y(N_FIFOCNT_1) );
    zao21b U1223 ( .A(_cell_531_U22_Z_0), .B(n3066), .C(n3194), .Y(n3088) );
    zmux21hb U1224 ( .A(TESTAD[3]), .B(TESTAD1135_3), .S(n2953), .Y(
        TESTAD1143_3) );
    zxo2b U1225 ( .A(add_362_carry_3), .B(TESTAD[3]), .Y(TESTAD1135_3) );
    zmux21hb U1226 ( .A(TESTAD[2]), .B(TESTAD1135_2), .S(n2953), .Y(
        TESTAD1143_2) );
    zhadrb add_362_U1_1_2 ( .A(TESTAD[2]), .B(add_362_carry_2), .CO(
        add_362_carry_3), .S(TESTAD1135_2) );
    zmux21hb U1227 ( .A(TESTAD[1]), .B(TESTAD1135_1), .S(n2953), .Y(
        TESTAD1143_1) );
    zhadrb add_362_U1_1_1 ( .A(TESTAD[1]), .B(TESTAD[0]), .CO(add_362_carry_2), 
        .S(TESTAD1135_1) );
    zmux21hb U1228 ( .A(ADI[31]), .B(PCIDATA_T_31), .S(n3215), .Y(
        PCIDATA_T1208_31) );
    zmux21hb U1229 ( .A(ADI[30]), .B(PCIDATA_T_30), .S(n3231), .Y(
        PCIDATA_T1208_30) );
    zmux21hb U1230 ( .A(ADI[29]), .B(PCIDATA_T_29), .S(n3215), .Y(
        PCIDATA_T1208_29) );
    zmux21hb U1231 ( .A(ADI[28]), .B(PCIDATA_T_28), .S(n3231), .Y(
        PCIDATA_T1208_28) );
    zmux21hb U1232 ( .A(ADI[27]), .B(PCIDATA_T_27), .S(n3215), .Y(
        PCIDATA_T1208_27) );
    zmux21hb U1233 ( .A(ADI[26]), .B(PCIDATA_T_26), .S(n3231), .Y(
        PCIDATA_T1208_26) );
    zmux21hb U1234 ( .A(ADI[25]), .B(PCIDATA_T_25), .S(n3215), .Y(
        PCIDATA_T1208_25) );
    zmux21hb U1235 ( .A(ADI[24]), .B(PCIDATA_T_24), .S(n3215), .Y(
        PCIDATA_T1208_24) );
    zmux21hb U1236 ( .A(ADI[23]), .B(PCIDATA_T_23), .S(n3231), .Y(
        PCIDATA_T1208_23) );
    zmux21hb U1237 ( .A(ADI[22]), .B(PCIDATA_T_22), .S(n3231), .Y(
        PCIDATA_T1208_22) );
    zmux21hb U1238 ( .A(ADI[21]), .B(PCIDATA_T_21), .S(n3215), .Y(
        PCIDATA_T1208_21) );
    zmux21hb U1239 ( .A(ADI[20]), .B(PCIDATA_T_20), .S(n3231), .Y(
        PCIDATA_T1208_20) );
    zmux21hb U1240 ( .A(ADI[19]), .B(PCIDATA_T_19), .S(n3215), .Y(
        PCIDATA_T1208_19) );
    zmux21hb U1241 ( .A(ADI[18]), .B(PCIDATA_T_18), .S(n3231), .Y(
        PCIDATA_T1208_18) );
    zmux21hb U1242 ( .A(ADI[17]), .B(PCIDATA_T_17), .S(n3231), .Y(
        PCIDATA_T1208_17) );
    zmux21hb U1243 ( .A(ADI[16]), .B(PCIDATA_T_16), .S(n3215), .Y(
        PCIDATA_T1208_16) );
    zmux21hb U1244 ( .A(ADI[15]), .B(PCIDATA_T_15), .S(n3231), .Y(
        PCIDATA_T1208_15) );
    zmux21hb U1245 ( .A(ADI[14]), .B(PCIDATA_T_14), .S(n3215), .Y(
        PCIDATA_T1208_14) );
    zmux21hb U1246 ( .A(ADI[13]), .B(PCIDATA_T_13), .S(n3231), .Y(
        PCIDATA_T1208_13) );
    zmux21hb U1247 ( .A(ADI[12]), .B(PCIDATA_T_12), .S(n3215), .Y(
        PCIDATA_T1208_12) );
    zmux21hb U1248 ( .A(ADI[11]), .B(PCIDATA_T_11), .S(n3231), .Y(
        PCIDATA_T1208_11) );
    zmux21hb U1249 ( .A(ADI[10]), .B(PCIDATA_T_10), .S(n3215), .Y(
        PCIDATA_T1208_10) );
    zmux21hb U1250 ( .A(ADI[9]), .B(PCIDATA_T_9), .S(n3231), .Y(
        PCIDATA_T1208_9) );
    zmux21hb U1251 ( .A(ADI[8]), .B(PCIDATA_T_8), .S(n3215), .Y(
        PCIDATA_T1208_8) );
    zmux21hb U1252 ( .A(ADI[7]), .B(PCIDATA_T_7), .S(n3231), .Y(
        PCIDATA_T1208_7) );
    zmux21hb U1253 ( .A(ADI[6]), .B(PCIDATA_T_6), .S(n3215), .Y(
        PCIDATA_T1208_6) );
    zmux21hb U1254 ( .A(ADI[5]), .B(PCIDATA_T_5), .S(n3231), .Y(
        PCIDATA_T1208_5) );
    zmux21hb U1255 ( .A(ADI[4]), .B(PCIDATA_T_4), .S(n3215), .Y(
        PCIDATA_T1208_4) );
    zmux21hb U1256 ( .A(ADI[3]), .B(PCIDATA_T_3), .S(n3231), .Y(
        PCIDATA_T1208_3) );
    zmux21hb U1257 ( .A(ADI[2]), .B(PCIDATA_T_2), .S(n3215), .Y(
        PCIDATA_T1208_2) );
    zmux21hb U1258 ( .A(ADI[1]), .B(PCIDATA_T_1), .S(n3231), .Y(
        PCIDATA_T1208_1) );
    zmux21hb U1259 ( .A(ADI[0]), .B(PCIDATA_T_0), .S(n3215), .Y(
        PCIDATA_T1208_0) );
    zao22b U1260 ( .A(rptr_8), .B(n3084), .C(c1328_9), .D(n2956), .Y(n_rptr_8)
         );
    zxo2b U1261 ( .A(add_416_carry_8), .B(rptr_8), .Y(c1328_9) );
    zao22b U1262 ( .A(rptr_7), .B(n3084), .C(c1328_8), .D(n2956), .Y(n_rptr_7)
         );
    zhadrb add_416_U1_1_7 ( .A(rptr_7), .B(add_416_carry_7), .CO(
        add_416_carry_8), .S(c1328_8) );
    zao22b U1263 ( .A(rptr_6), .B(n3084), .C(c1328_7), .D(n2956), .Y(n_rptr_6)
         );
    zhadrb add_416_U1_1_6 ( .A(rptr_6), .B(add_416_carry_6), .CO(
        add_416_carry_7), .S(c1328_7) );
    zao22b U1264 ( .A(rptr_5), .B(n3084), .C(c1328_6), .D(n2956), .Y(n_rptr_5)
         );
    zhadrb add_416_U1_1_5 ( .A(rptr_5), .B(add_416_carry_5), .CO(
        add_416_carry_6), .S(c1328_6) );
    zao22b U1265 ( .A(rptr_4), .B(n3084), .C(c1328_5), .D(n2956), .Y(n_rptr_4)
         );
    zhadrb add_416_U1_1_4 ( .A(rptr_4), .B(add_416_carry_4), .CO(
        add_416_carry_5), .S(c1328_5) );
    zao22b U1266 ( .A(rptr_3), .B(n3084), .C(c1328_4), .D(n2956), .Y(n_rptr_3)
         );
    zhadrb add_416_U1_1_3 ( .A(rptr_3), .B(add_416_carry_3), .CO(
        add_416_carry_4), .S(c1328_4) );
    zao22b U1267 ( .A(rptr_2), .B(n3084), .C(c1328_3), .D(n2956), .Y(n_rptr_2)
         );
    zhadrb add_416_U1_1_2 ( .A(rptr_2), .B(add_416_carry_2), .CO(
        add_416_carry_3), .S(c1328_3) );
    zao22b U1268 ( .A(rptr_0), .B(n3084), .C(c1328_1), .D(n2956), .Y(n_rptr_0)
         );
    zor2b U1269 ( .A(n3085), .B(n3066), .Y(n3084) );
    zao22b U1270 ( .A(FSIZE_1), .B(n2954), .C(FSIZE1554_1), .D(n3087), .Y(
        FSIZE1570_1) );
    zxo3b r255_U1_1 ( .A(FSIZE_1), .B(_cell_531_U41_Z_0), .C(r255_carry_1), 
        .Y(FSIZE1554_1) );
    zao22b U1271 ( .A(FSIZE_0), .B(n2954), .C(FSIZE1554_0), .D(n3087), .Y(
        FSIZE1570_0) );
    zor2b U1272 ( .A(n3001), .B(n3199), .Y(n3087) );
    zmux21hb U1273 ( .A(MDO[31]), .B(FFRDPCI[31]), .S(n3217), .Y(
        FFRDPCI1761_31) );
    zmux21hb U1274 ( .A(MDO[30]), .B(FFRDPCI[30]), .S(n3225), .Y(
        FFRDPCI1761_30) );
    zmux21hb U1275 ( .A(MDO[29]), .B(FFRDPCI[29]), .S(n3217), .Y(
        FFRDPCI1761_29) );
    zmux21hb U1276 ( .A(MDO[28]), .B(FFRDPCI[28]), .S(n3225), .Y(
        FFRDPCI1761_28) );
    zmux21hb U1277 ( .A(MDO[27]), .B(FFRDPCI[27]), .S(n3217), .Y(
        FFRDPCI1761_27) );
    zmux21hb U1278 ( .A(MDO[26]), .B(FFRDPCI[26]), .S(n3225), .Y(
        FFRDPCI1761_26) );
    zmux21hb U1279 ( .A(MDO[25]), .B(FFRDPCI[25]), .S(n3217), .Y(
        FFRDPCI1761_25) );
    zmux21hb U1280 ( .A(MDO[24]), .B(FFRDPCI[24]), .S(n3217), .Y(
        FFRDPCI1761_24) );
    zmux21hb U1281 ( .A(MDO[23]), .B(FFRDPCI[23]), .S(n3225), .Y(
        FFRDPCI1761_23) );
    zmux21hb U1282 ( .A(MDO[22]), .B(FFRDPCI[22]), .S(n3225), .Y(
        FFRDPCI1761_22) );
    zmux21hb U1283 ( .A(MDO[21]), .B(FFRDPCI[21]), .S(n3217), .Y(
        FFRDPCI1761_21) );
    zmux21hb U1284 ( .A(MDO[20]), .B(FFRDPCI[20]), .S(n3225), .Y(
        FFRDPCI1761_20) );
    zmux21hb U1285 ( .A(MDO[19]), .B(FFRDPCI[19]), .S(n3217), .Y(
        FFRDPCI1761_19) );
    zmux21hb U1286 ( .A(MDO[18]), .B(FFRDPCI[18]), .S(n3225), .Y(
        FFRDPCI1761_18) );
    zmux21hb U1287 ( .A(MDO[17]), .B(FFRDPCI[17]), .S(n3225), .Y(
        FFRDPCI1761_17) );
    zmux21hb U1288 ( .A(MDO[16]), .B(FFRDPCI[16]), .S(n3217), .Y(
        FFRDPCI1761_16) );
    zmux21hb U1289 ( .A(MDO[15]), .B(FFRDPCI[15]), .S(n3225), .Y(
        FFRDPCI1761_15) );
    zmux21hb U1290 ( .A(MDO[14]), .B(FFRDPCI[14]), .S(n3217), .Y(
        FFRDPCI1761_14) );
    zmux21hb U1291 ( .A(MDO[13]), .B(FFRDPCI[13]), .S(n3225), .Y(
        FFRDPCI1761_13) );
    zmux21hb U1292 ( .A(MDO[12]), .B(FFRDPCI[12]), .S(n3217), .Y(
        FFRDPCI1761_12) );
    zmux21hb U1293 ( .A(MDO[11]), .B(FFRDPCI[11]), .S(n3225), .Y(
        FFRDPCI1761_11) );
    zmux21hb U1294 ( .A(MDO[10]), .B(FFRDPCI[10]), .S(n3217), .Y(
        FFRDPCI1761_10) );
    zmux21hb U1295 ( .A(MDO[9]), .B(FFRDPCI[9]), .S(n3225), .Y(FFRDPCI1761_9)
         );
    zmux21hb U1296 ( .A(MDO[8]), .B(FFRDPCI[8]), .S(n3217), .Y(FFRDPCI1761_8)
         );
    zmux21hb U1297 ( .A(MDO[7]), .B(FFRDPCI[7]), .S(n3225), .Y(FFRDPCI1761_7)
         );
    zmux21hb U1298 ( .A(MDO[6]), .B(FFRDPCI[6]), .S(n3217), .Y(FFRDPCI1761_6)
         );
    zmux21hb U1299 ( .A(MDO[5]), .B(FFRDPCI[5]), .S(n3225), .Y(FFRDPCI1761_5)
         );
    zmux21hb U1300 ( .A(MDO[4]), .B(FFRDPCI[4]), .S(n3217), .Y(FFRDPCI1761_4)
         );
    zmux21hb U1301 ( .A(MDO[3]), .B(FFRDPCI[3]), .S(n3225), .Y(FFRDPCI1761_3)
         );
    zmux21hb U1302 ( .A(MDO[2]), .B(FFRDPCI[2]), .S(n3217), .Y(FFRDPCI1761_2)
         );
    zmux21hb U1303 ( .A(MDO[1]), .B(FFRDPCI[1]), .S(n3225), .Y(FFRDPCI1761_1)
         );
    zmux21hb U1304 ( .A(MDO[0]), .B(FFRDPCI[0]), .S(n3217), .Y(FFRDPCI1761_0)
         );
    zivb U1305 ( .A(n3224), .Y(n3217) );
    zor2b U1306 ( .A(PCIREAD), .B(n2949), .Y(n3224) );
    zivb U1307 ( .A(n3224), .Y(n3225) );
    zmux21lb U1308 ( .A(n3189), .B(n3208), .S(n2998), .Y(TCNT1958_1) );
    zmux21lb U1309 ( .A(n2587), .B(TCNT1929_1), .S(UPOP), .Y(n3208) );
    zmux21lb U1310 ( .A(n3189), .B(n3210), .S(LDWPR), .Y(ST_BE2037_1) );
    zivb U1311 ( .A(WPR1), .Y(n3210) );
    zmux21lb U1312 ( .A(n3191), .B(n3211), .S(LDWPR), .Y(ST_BE2037_0) );
    zivb U1313 ( .A(WPR0), .Y(n3211) );
    zivb U1314 ( .A(n3110), .Y(n3077) );
    zor2b U1315 ( .A(RCNT_1), .B(n3102), .Y(n3110) );
    zao22b U1316 ( .A(UCBEO_[0]), .B(n2951), .C(n2958), .D(END_BE_0), .Y(
        END_BE2076_0) );
    zivb U1317 ( .A(PCIWRT), .Y(n3206) );
    zmux21hb U1318 ( .A(MDO[31]), .B(FFRDUSB_31), .S(n3216), .Y(FFRDUSB2141_31
        ) );
    zmux21hb U1319 ( .A(MDO[30]), .B(FFRDUSB_30), .S(n3226), .Y(FFRDUSB2141_30
        ) );
    zmux21hb U1320 ( .A(MDO[29]), .B(FFRDUSB_29), .S(n3216), .Y(FFRDUSB2141_29
        ) );
    zmux21hb U1321 ( .A(MDO[28]), .B(FFRDUSB_28), .S(n3226), .Y(FFRDUSB2141_28
        ) );
    zmux21hb U1322 ( .A(MDO[27]), .B(FFRDUSB_27), .S(n3216), .Y(FFRDUSB2141_27
        ) );
    zmux21hb U1323 ( .A(MDO[26]), .B(FFRDUSB_26), .S(n3226), .Y(FFRDUSB2141_26
        ) );
    zmux21hb U1324 ( .A(MDO[25]), .B(FFRDUSB_25), .S(n3216), .Y(FFRDUSB2141_25
        ) );
    zmux21hb U1325 ( .A(MDO[24]), .B(FFRDUSB_24), .S(n3226), .Y(FFRDUSB2141_24
        ) );
    zmux21hb U1326 ( .A(MDO[23]), .B(FFRDUSB_23), .S(n3216), .Y(FFRDUSB2141_23
        ) );
    zmux21hb U1327 ( .A(MDO[22]), .B(FFRDUSB_22), .S(n3226), .Y(FFRDUSB2141_22
        ) );
    zmux21hb U1328 ( .A(MDO[21]), .B(FFRDUSB_21), .S(n3216), .Y(FFRDUSB2141_21
        ) );
    zmux21hb U1329 ( .A(MDO[20]), .B(FFRDUSB_20), .S(n3226), .Y(FFRDUSB2141_20
        ) );
    zmux21hb U1330 ( .A(MDO[19]), .B(FFRDUSB_19), .S(n3226), .Y(FFRDUSB2141_19
        ) );
    zmux21hb U1331 ( .A(MDO[18]), .B(FFRDUSB_18), .S(n3216), .Y(FFRDUSB2141_18
        ) );
    zmux21hb U1332 ( .A(MDO[17]), .B(FFRDUSB_17), .S(n3226), .Y(FFRDUSB2141_17
        ) );
    zmux21hb U1333 ( .A(MDO[16]), .B(FFRDUSB_16), .S(n3216), .Y(FFRDUSB2141_16
        ) );
    zmux21hb U1334 ( .A(MDO[15]), .B(FFRDUSB_15), .S(n3226), .Y(FFRDUSB2141_15
        ) );
    zmux21hb U1335 ( .A(MDO[14]), .B(FFRDUSB_14), .S(n3216), .Y(FFRDUSB2141_14
        ) );
    zmux21hb U1336 ( .A(MDO[13]), .B(FFRDUSB_13), .S(n3226), .Y(FFRDUSB2141_13
        ) );
    zmux21hb U1337 ( .A(MDO[12]), .B(FFRDUSB_12), .S(n3216), .Y(FFRDUSB2141_12
        ) );
    zmux21hb U1338 ( .A(MDO[11]), .B(FFRDUSB_11), .S(n3216), .Y(FFRDUSB2141_11
        ) );
    zmux21hb U1339 ( .A(MDO[10]), .B(FFRDUSB_10), .S(n3226), .Y(FFRDUSB2141_10
        ) );
    zmux21hb U1340 ( .A(MDO[9]), .B(FFRDUSB_9), .S(n3226), .Y(FFRDUSB2141_9)
         );
    zmux21hb U1341 ( .A(MDO[8]), .B(FFRDUSB_8), .S(n3216), .Y(FFRDUSB2141_8)
         );
    zmux21hb U1342 ( .A(MDO[7]), .B(FFRDUSB_7), .S(n3226), .Y(FFRDUSB2141_7)
         );
    zmux21hb U1343 ( .A(MDO[6]), .B(FFRDUSB_6), .S(n3216), .Y(FFRDUSB2141_6)
         );
    zmux21hb U1344 ( .A(MDO[5]), .B(FFRDUSB_5), .S(n3226), .Y(FFRDUSB2141_5)
         );
    zmux21hb U1345 ( .A(MDO[4]), .B(FFRDUSB_4), .S(n3216), .Y(FFRDUSB2141_4)
         );
    zmux21hb U1346 ( .A(MDO[3]), .B(FFRDUSB_3), .S(n3226), .Y(FFRDUSB2141_3)
         );
    zmux21hb U1347 ( .A(MDO[2]), .B(FFRDUSB_2), .S(n3216), .Y(FFRDUSB2141_2)
         );
    zmux21hb U1348 ( .A(MDO[1]), .B(FFRDUSB_1), .S(n3216), .Y(FFRDUSB2141_1)
         );
    zmux21hb U1349 ( .A(MDO[0]), .B(FFRDUSB_0), .S(n3226), .Y(FFRDUSB2141_0)
         );
    zivb U1350 ( .A(n3223), .Y(n3226) );
    zivb U1351 ( .A(n3223), .Y(n3216) );
    zor2b U1352 ( .A(FEMPTY), .B(n3203), .Y(n3071) );
    zivb U1353 ( .A(n3071), .Y(n3202) );
    zan2b U1354 ( .A(END_BE_1), .B(n3071), .Y(n3070) );
    zor2b U1355 ( .A(PROCESS), .B(n3006), .Y(PROCESS2334) );
    zivb U1356 ( .A(n3186), .Y(PCIWRT_TEST1184) );
    zivb U1357 ( .A(n3021), .Y(n3029) );
    zao21b U1358 ( .A(USBREAD), .B(n3066), .C(n3067), .Y(FPOP_T1737) );
    zao21b U1359 ( .A(RDFFNXT_1), .B(n3068), .C(n2960), .Y(n3067) );
    zivb U1360 ( .A(n3067), .Y(n3086) );
    zao32b U1361 ( .A(PROCESS), .B(n3064), .C(n3000), .D(EOT3_T), .E(FEMPTY), 
        .Y(EOT3_T1447) );
    zivb U1362 ( .A(EOT), .Y(n3193) );
    zmux21lb U1363 ( .A(n3091), .B(n3212), .S(n3090), .Y(RXPKTEND_T2371) );
    zor2b U1364 ( .A(RXPKTEND), .B(n3083), .Y(n3212) );
    znr2b U1365 ( .A(RXERR), .B(EOT), .Y(n3090) );
    zoai21b U1366 ( .A(RDMAEND), .B(n3082), .C(n3083), .Y(RXPKTEND2408) );
    zivb U1367 ( .A(n3021), .Y(n3028) );
    zivb U1368 ( .A(n3103), .Y(n3075) );
    zor2b U1369 ( .A(n3101), .B(n3102), .Y(n3103) );
    zor2b U1370 ( .A(FPOP), .B(FPOP_ONCE), .Y(FPOP_ONCE1612) );
    zivb U1371 ( .A(n3021), .Y(n3030) );
    zor2b U1372 ( .A(PCIWRT_TEST), .B(PCIWRT), .Y(PSH1244) );
    zivb U1373 ( .A(PSH1244), .Y(n3215) );
    zivb U1374 ( .A(PSH1244), .Y(n3231) );
    zivb U1375 ( .A(n3021), .Y(n3031) );
    zivb U1376 ( .A(n3021), .Y(n3027) );
    zan2b U1377 ( .A(PROCESS), .B(n3064), .Y(n3096) );
    zivb U1378 ( .A(n3105), .Y(n3085) );
    zor2b U1379 ( .A(FIFOCNT_1), .B(n3097), .Y(n3098) );
    zivb U1380 ( .A(n3196), .Y(n3227) );
    zor2b U1381 ( .A(RXFIFO), .B(n3228), .Y(n3196) );
    zivb U1382 ( .A(n3003), .Y(n3228) );
    zivb U1383 ( .A(n3003), .Y(n3229) );
    zivb U1384 ( .A(n3197), .Y(n3081) );
    zor2b U1385 ( .A(n3004), .B(n3100), .Y(n3197) );
    zivb U1386 ( .A(RXFIFO), .Y(n3100) );
    zivb U1387 ( .A(n3196), .Y(n3080) );
    zivb U1388 ( .A(n3197), .Y(n3230) );
    zor2b U1389 ( .A(PCIREAD), .B(FPOP_T), .Y(FPOP) );
    zivb U1390 ( .A(FPOP), .Y(n3066) );
    zmux41b U1391 ( .A(n2586), .B(n2587), .D0(FFRDUSB_0), .D1(FFRDUSB_8), .D2(
        FFRDUSB_16), .D3(FFRDUSB_24), .Y(HOSTDAT[0]) );
    zmux41b U1392 ( .A(n2586), .B(n2587), .D0(FFRDUSB_1), .D1(FFRDUSB_9), .D2(
        FFRDUSB_17), .D3(FFRDUSB_25), .Y(HOSTDAT[1]) );
    zmux41b U1393 ( .A(n2586), .B(n2587), .D0(FFRDUSB_2), .D1(FFRDUSB_10), 
        .D2(FFRDUSB_18), .D3(FFRDUSB_26), .Y(HOSTDAT[2]) );
    zmux41b U1394 ( .A(n2586), .B(n2587), .D0(FFRDUSB_3), .D1(FFRDUSB_11), 
        .D2(FFRDUSB_19), .D3(FFRDUSB_27), .Y(HOSTDAT[3]) );
    zmux41b U1395 ( .A(n2586), .B(n2587), .D0(FFRDUSB_4), .D1(FFRDUSB_12), 
        .D2(FFRDUSB_20), .D3(FFRDUSB_28), .Y(HOSTDAT[4]) );
    zmux41b U1396 ( .A(n2586), .B(n2587), .D0(FFRDUSB_5), .D1(FFRDUSB_13), 
        .D2(FFRDUSB_21), .D3(FFRDUSB_29), .Y(HOSTDAT[5]) );
    zmux41b U1397 ( .A(n2586), .B(n2587), .D0(FFRDUSB_6), .D1(FFRDUSB_14), 
        .D2(FFRDUSB_22), .D3(FFRDUSB_30), .Y(HOSTDAT[6]) );
    zmux41b U1398 ( .A(n2586), .B(n2587), .D0(FFRDUSB_7), .D1(FFRDUSB_15), 
        .D2(FFRDUSB_23), .D3(FFRDUSB_31), .Y(HOSTDAT[7]) );
    zivb U1399 ( .A(FIFOCNT_0), .Y(n3093) );
    zivb U1400 ( .A(USBFFTMP_6), .Y(n3154) );
    zivb U1401 ( .A(USBFFTMP_25), .Y(n3164) );
    zivb U1402 ( .A(USBFFTMP_15), .Y(n3175) );
    zivb U1403 ( .A(USBFFTMP_26), .Y(n3163) );
    zivb U1404 ( .A(FIFO_OK), .Y(n3074) );
    zivb U1405 ( .A(USBFFTMP_19), .Y(n3171) );
    zivb U1406 ( .A(USBFFTMP_21), .Y(n3168) );
    zivb U1407 ( .A(USBFFTMP_14), .Y(n3176) );
    zivb U1408 ( .A(USBFFTMP_30), .Y(n3158) );
    zivb U1409 ( .A(USBFFTMP_10), .Y(n3180) );
    zdffqrb RCNT_reg_1 ( .CK(CLK60M), .D(RCNT351_1), .R(n3028), .Q(RCNT_1) );
    zivb U1410 ( .A(RCNT_1), .Y(n3101) );
    zdffrb USBTMP_reg_31 ( .CK(CLK60M), .D(USBTMP396_31), .R(n3028), .QN(n3122
        ) );
    zdffrb USBTMP_reg_29 ( .CK(CLK60M), .D(USBTMP396_29), .R(n3024), .QN(n3126
        ) );
    zdffrb USBTMP_reg_28 ( .CK(CLK60M), .D(USBTMP396_28), .R(n3030), .QN(n3127
        ) );
    zdffrb USBTMP_reg_27 ( .CK(CLK60M), .D(USBTMP396_27), .R(n3030), .QN(n3128
        ) );
    zdffrb USBTMP_reg_26 ( .CK(CLK60M), .D(USBTMP396_26), .R(n3023), .QN(n3129
        ) );
    zdffrb USBTMP_reg_25 ( .CK(CLK60M), .D(USBTMP396_25), .R(n3027), .QN(n3131
        ) );
    zdffrb USBTMP_reg_23 ( .CK(CLK60M), .D(USBTMP396_23), .R(n3026), .QN(n3133
        ) );
    zdffrb USBTMP_reg_22 ( .CK(CLK60M), .D(USBTMP396_22), .R(n3024), .QN(n3135
        ) );
    zdffrb USBTMP_reg_21 ( .CK(CLK60M), .D(USBTMP396_21), .R(n3026), .QN(n3136
        ) );
    zdffrb USBTMP_reg_20 ( .CK(CLK60M), .D(USBTMP396_20), .R(n3025), .QN(n3137
        ) );
    zdffrb USBTMP_reg_19 ( .CK(CLK60M), .D(USBTMP396_19), .R(n3028), .QN(n3139
        ) );
    zdffrb USBTMP_reg_18 ( .CK(CLK60M), .D(USBTMP396_18), .R(n3026), .QN(n3140
        ) );
    zdffrb USBTMP_reg_17 ( .CK(CLK60M), .D(USBTMP396_17), .R(n3022), .QN(n3141
        ) );
    zdffrb USBTMP_reg_15 ( .CK(CLK60M), .D(USBTMP396_15), .R(n3029), .QN(n3143
        ) );
    zdffrb USBTMP_reg_14 ( .CK(CLK60M), .D(USBTMP396_14), .R(n3024), .QN(n3144
        ) );
    zdffrb USBTMP_reg_10 ( .CK(CLK60M), .D(USBTMP396_10), .R(n3029), .QN(n3148
        ) );
    zdffrb USBTMP_reg_8 ( .CK(CLK60M), .D(USBTMP396_8), .R(n3031), .QN(n3111)
         );
    zdffrb USBTMP_reg_6 ( .CK(CLK60M), .D(USBTMP396_6), .R(n3027), .QN(n3116)
         );
    zdffrb USBTMP_reg_5 ( .CK(CLK60M), .D(USBTMP396_5), .R(n3022), .QN(n3118)
         );
    zdffrb USBTMP_reg_4 ( .CK(CLK60M), .D(USBTMP396_4), .R(n3029), .QN(n3120)
         );
    zdffrb USBTMP_reg_3 ( .CK(CLK60M), .D(USBTMP396_3), .R(n3031), .QN(n3124)
         );
    zdffrb USBTMP_reg_2 ( .CK(CLK60M), .D(USBTMP396_2), .R(n3023), .QN(n3138)
         );
    zdffrb USBTMP_reg_1 ( .CK(CLK60M), .D(USBTMP396_1), .R(n3028), .QN(n3149)
         );
    zdffqrb USBFFTMP_reg_31 ( .CK(CLK60M), .D(USBFFTMP655_31), .R(n3028), .Q(
        USBFFTMP_31) );
    zivb U1411 ( .A(USBFFTMP_31), .Y(n3157) );
    zdffqrb USBFFTMP_reg_29 ( .CK(CLK60M), .D(USBFFTMP655_29), .R(n3023), .Q(
        USBFFTMP_29) );
    zivb U1412 ( .A(USBFFTMP_29), .Y(n3160) );
    zdffqrb USBFFTMP_reg_28 ( .CK(CLK60M), .D(USBFFTMP655_28), .R(n3026), .Q(
        USBFFTMP_28) );
    zivb U1413 ( .A(USBFFTMP_28), .Y(n3161) );
    zdffqrb USBFFTMP_reg_27 ( .CK(CLK60M), .D(USBFFTMP655_27), .R(n3025), .Q(
        USBFFTMP_27) );
    zivb U1414 ( .A(USBFFTMP_27), .Y(n3162) );
    zdffqrb USBFFTMP_reg_24 ( .CK(CLK60M), .D(USBFFTMP655_24), .R(n3023), .Q(
        USBFFTMP_24) );
    zivb U1415 ( .A(USBFFTMP_24), .Y(n3165) );
    zdffqrb USBFFTMP_reg_23 ( .CK(CLK60M), .D(USBFFTMP655_23), .R(n3023), .Q(
        USBFFTMP_23) );
    zivb U1416 ( .A(USBFFTMP_23), .Y(n3166) );
    zdffqrb USBFFTMP_reg_22 ( .CK(CLK60M), .D(USBFFTMP655_22), .R(n3031), .Q(
        USBFFTMP_22) );
    zivb U1417 ( .A(USBFFTMP_22), .Y(n3167) );
    zdffqrb USBFFTMP_reg_20 ( .CK(CLK60M), .D(USBFFTMP655_20), .R(n3027), .Q(
        USBFFTMP_20) );
    zivb U1418 ( .A(USBFFTMP_20), .Y(n3169) );
    zdffqrb USBFFTMP_reg_18 ( .CK(CLK60M), .D(USBFFTMP655_18), .R(n3024), .Q(
        USBFFTMP_18) );
    zivb U1419 ( .A(USBFFTMP_18), .Y(n3172) );
    zdffqrb USBFFTMP_reg_17 ( .CK(CLK60M), .D(USBFFTMP655_17), .R(n3024), .Q(
        USBFFTMP_17) );
    zivb U1420 ( .A(USBFFTMP_17), .Y(n3173) );
    zdffqrb USBFFTMP_reg_16 ( .CK(CLK60M), .D(USBFFTMP655_16), .R(n3030), .Q(
        USBFFTMP_16) );
    zivb U1421 ( .A(USBFFTMP_16), .Y(n3174) );
    zdffqrb USBFFTMP_reg_13 ( .CK(CLK60M), .D(USBFFTMP655_13), .R(n3025), .Q(
        USBFFTMP_13) );
    zivb U1422 ( .A(USBFFTMP_13), .Y(n3177) );
    zdffqrb USBFFTMP_reg_12 ( .CK(CLK60M), .D(USBFFTMP655_12), .R(n3022), .Q(
        USBFFTMP_12) );
    zivb U1423 ( .A(USBFFTMP_12), .Y(n3178) );
    zdffqrb USBFFTMP_reg_11 ( .CK(CLK60M), .D(USBFFTMP655_11), .R(n3027), .Q(
        USBFFTMP_11) );
    zivb U1424 ( .A(USBFFTMP_11), .Y(n3179) );
    zdffqrb USBFFTMP_reg_9 ( .CK(CLK60M), .D(USBFFTMP655_9), .R(n3022), .Q(
        USBFFTMP_9) );
    zivb U1425 ( .A(USBFFTMP_9), .Y(n3151) );
    zdffqrb USBFFTMP_reg_8 ( .CK(CLK60M), .D(USBFFTMP655_8), .R(n3024), .Q(
        USBFFTMP_8) );
    zivb U1426 ( .A(USBFFTMP_8), .Y(n3152) );
    zdffqrb USBFFTMP_reg_7 ( .CK(CLK60M), .D(USBFFTMP655_7), .R(n3030), .Q(
        USBFFTMP_7) );
    zivb U1427 ( .A(USBFFTMP_7), .Y(n3153) );
    zdffqrb USBFFTMP_reg_5 ( .CK(CLK60M), .D(USBFFTMP655_5), .R(n3029), .Q(
        USBFFTMP_5) );
    zivb U1428 ( .A(USBFFTMP_5), .Y(n3155) );
    zdffqrb USBFFTMP_reg_4 ( .CK(CLK60M), .D(USBFFTMP655_4), .R(n3022), .Q(
        USBFFTMP_4) );
    zivb U1429 ( .A(USBFFTMP_4), .Y(n3156) );
    zdffqrb USBFFTMP_reg_3 ( .CK(CLK60M), .D(USBFFTMP655_3), .R(n3028), .Q(
        USBFFTMP_3) );
    zivb U1430 ( .A(USBFFTMP_3), .Y(n3159) );
    zdffqrb USBFFTMP_reg_2 ( .CK(CLK60M), .D(USBFFTMP655_2), .R(n3031), .Q(
        USBFFTMP_2) );
    zivb U1431 ( .A(USBFFTMP_2), .Y(n3170) );
    zdffqrb USBFFTMP_reg_1 ( .CK(CLK60M), .D(USBFFTMP655_1), .R(n3025), .Q(
        USBFFTMP_1) );
    zivb U1432 ( .A(USBFFTMP_1), .Y(n3181) );
    zdffqrb USBFFTMP_reg_0 ( .CK(CLK60M), .D(USBFFTMP655_0), .R(n3029), .Q(
        USBFFTMP_0) );
    zivb U1433 ( .A(USBFFTMP_0), .Y(n3182) );
    zdffqrb FIFOCNT_reg_8 ( .CK(PCICLK), .D(N_FIFOCNT_8), .R(n3026), .Q(
        FIFOCNT_8) );
    zivb U1434 ( .A(FIFOCNT_8), .Y(n3094) );
    zdffqrb FIFOCNT_reg_7 ( .CK(PCICLK), .D(N_FIFOCNT_7), .R(n3023), .Q(
        FIFOCNT_7) );
    zdffqrb FIFOCNT_reg_6 ( .CK(PCICLK), .D(N_FIFOCNT_6), .R(n3026), .Q(
        FIFOCNT_6) );
    zdffqrb FIFOCNT_reg_5 ( .CK(PCICLK), .D(N_FIFOCNT_5), .R(n3023), .Q(
        FIFOCNT_5) );
    zdffqrb FIFOCNT_reg_4 ( .CK(PCICLK), .D(N_FIFOCNT_4), .R(n3026), .Q(
        FIFOCNT_4) );
    zdffqrb FIFOCNT_reg_3 ( .CK(PCICLK), .D(N_FIFOCNT_3), .R(n3025), .Q(
        FIFOCNT_3) );
    zdffqrb FIFOCNT_reg_2 ( .CK(PCICLK), .D(N_FIFOCNT_2), .R(n3023), .Q(
        FIFOCNT_2) );
    zdffqrb FIFOCNT_reg_1 ( .CK(PCICLK), .D(N_FIFOCNT_1), .R(n3030), .Q(
        FIFOCNT_1) );
    zdffqrb_ WMA_reg_6 ( .CK(PCICLK), .D(wptr_6), .R(n3022), .Q(WMA[6]) );
    zdffqrb_ WMA_reg_4 ( .CK(PCICLK), .D(wptr_4), .R(n3030), .Q(WMA[4]) );
    zdffqrb_ WMA_reg_3 ( .CK(PCICLK), .D(wptr_3), .R(n3031), .Q(WMA[3]) );
    zdffqrb_ WMA_reg_2 ( .CK(PCICLK), .D(wptr_2), .R(n3027), .Q(WMA[2]) );
    zdffqrb_ WMA_reg_1 ( .CK(PCICLK), .D(wptr_1), .R(n3029), .Q(WMA[1]) );
    zdffqrb_ WMA_reg_0 ( .CK(PCICLK), .D(wptr_0), .R(n3027), .Q(WMA[0]) );
    zdffqrb TESTAD_reg_3 ( .CK(PCICLK), .D(TESTAD1143_3), .R(n3007), .Q(TESTAD
        [3]) );
    zivb U1435 ( .A(TESTAD[3]), .Y(n3184) );
    zdffqrb TESTAD_reg_2 ( .CK(PCICLK), .D(TESTAD1143_2), .R(n3007), .Q(TESTAD
        [2]) );
    zivb U1436 ( .A(TESTAD[2]), .Y(n3185) );
    zdffqrb TESTAD_reg_1 ( .CK(PCICLK), .D(TESTAD1143_1), .R(n3007), .Q(TESTAD
        [1]) );
    zdffqb PCIDATA_T_reg_31 ( .CK(PCICLK), .D(PCIDATA_T1208_31), .Q(
        PCIDATA_T_31) );
    zdffqb PCIDATA_T_reg_30 ( .CK(PCICLK), .D(PCIDATA_T1208_30), .Q(
        PCIDATA_T_30) );
    zdffqb PCIDATA_T_reg_29 ( .CK(PCICLK), .D(PCIDATA_T1208_29), .Q(
        PCIDATA_T_29) );
    zdffqb PCIDATA_T_reg_28 ( .CK(PCICLK), .D(PCIDATA_T1208_28), .Q(
        PCIDATA_T_28) );
    zdffqb PCIDATA_T_reg_27 ( .CK(PCICLK), .D(PCIDATA_T1208_27), .Q(
        PCIDATA_T_27) );
    zdffqb PCIDATA_T_reg_26 ( .CK(PCICLK), .D(PCIDATA_T1208_26), .Q(
        PCIDATA_T_26) );
    zdffqb PCIDATA_T_reg_25 ( .CK(PCICLK), .D(PCIDATA_T1208_25), .Q(
        PCIDATA_T_25) );
    zdffqb PCIDATA_T_reg_24 ( .CK(PCICLK), .D(PCIDATA_T1208_24), .Q(
        PCIDATA_T_24) );
    zdffqb PCIDATA_T_reg_23 ( .CK(PCICLK), .D(PCIDATA_T1208_23), .Q(
        PCIDATA_T_23) );
    zdffqb PCIDATA_T_reg_22 ( .CK(PCICLK), .D(PCIDATA_T1208_22), .Q(
        PCIDATA_T_22) );
    zdffqb PCIDATA_T_reg_21 ( .CK(PCICLK), .D(PCIDATA_T1208_21), .Q(
        PCIDATA_T_21) );
    zdffqb PCIDATA_T_reg_20 ( .CK(PCICLK), .D(PCIDATA_T1208_20), .Q(
        PCIDATA_T_20) );
    zdffqb PCIDATA_T_reg_19 ( .CK(PCICLK), .D(PCIDATA_T1208_19), .Q(
        PCIDATA_T_19) );
    zdffqb PCIDATA_T_reg_18 ( .CK(PCICLK), .D(PCIDATA_T1208_18), .Q(
        PCIDATA_T_18) );
    zdffqb PCIDATA_T_reg_17 ( .CK(PCICLK), .D(PCIDATA_T1208_17), .Q(
        PCIDATA_T_17) );
    zdffqb PCIDATA_T_reg_16 ( .CK(PCICLK), .D(PCIDATA_T1208_16), .Q(
        PCIDATA_T_16) );
    zdffqb PCIDATA_T_reg_15 ( .CK(PCICLK), .D(PCIDATA_T1208_15), .Q(
        PCIDATA_T_15) );
    zdffqb PCIDATA_T_reg_14 ( .CK(PCICLK), .D(PCIDATA_T1208_14), .Q(
        PCIDATA_T_14) );
    zdffqb PCIDATA_T_reg_13 ( .CK(PCICLK), .D(PCIDATA_T1208_13), .Q(
        PCIDATA_T_13) );
    zdffqb PCIDATA_T_reg_12 ( .CK(PCICLK), .D(PCIDATA_T1208_12), .Q(
        PCIDATA_T_12) );
    zdffqb PCIDATA_T_reg_11 ( .CK(PCICLK), .D(PCIDATA_T1208_11), .Q(
        PCIDATA_T_11) );
    zdffqb PCIDATA_T_reg_10 ( .CK(PCICLK), .D(PCIDATA_T1208_10), .Q(
        PCIDATA_T_10) );
    zdffqb PCIDATA_T_reg_9 ( .CK(PCICLK), .D(PCIDATA_T1208_9), .Q(PCIDATA_T_9)
         );
    zdffqb PCIDATA_T_reg_8 ( .CK(PCICLK), .D(PCIDATA_T1208_8), .Q(PCIDATA_T_8)
         );
    zdffqb PCIDATA_T_reg_7 ( .CK(PCICLK), .D(PCIDATA_T1208_7), .Q(PCIDATA_T_7)
         );
    zdffqb PCIDATA_T_reg_6 ( .CK(PCICLK), .D(PCIDATA_T1208_6), .Q(PCIDATA_T_6)
         );
    zdffqb PCIDATA_T_reg_5 ( .CK(PCICLK), .D(PCIDATA_T1208_5), .Q(PCIDATA_T_5)
         );
    zdffqb PCIDATA_T_reg_4 ( .CK(PCICLK), .D(PCIDATA_T1208_4), .Q(PCIDATA_T_4)
         );
    zdffqb PCIDATA_T_reg_3 ( .CK(PCICLK), .D(PCIDATA_T1208_3), .Q(PCIDATA_T_3)
         );
    zdffqb PCIDATA_T_reg_2 ( .CK(PCICLK), .D(PCIDATA_T1208_2), .Q(PCIDATA_T_2)
         );
    zdffqb PCIDATA_T_reg_1 ( .CK(PCICLK), .D(PCIDATA_T1208_1), .Q(PCIDATA_T_1)
         );
    zdffqb PCIDATA_T_reg_0 ( .CK(PCICLK), .D(PCIDATA_T1208_0), .Q(PCIDATA_T_0)
         );
    zdffqb_ PCIDATA_reg_31 ( .CK(PCICLK), .D(PCIDATA_T_31), .Q(PCIDATA_31) );
    zdffqb_ PCIDATA_reg_30 ( .CK(PCICLK), .D(PCIDATA_T_30), .Q(PCIDATA_30) );
    zdffqb_ PCIDATA_reg_29 ( .CK(PCICLK), .D(PCIDATA_T_29), .Q(PCIDATA_29) );
    zdffqb_ PCIDATA_reg_28 ( .CK(PCICLK), .D(PCIDATA_T_28), .Q(PCIDATA_28) );
    zdffqb_ PCIDATA_reg_27 ( .CK(PCICLK), .D(PCIDATA_T_27), .Q(PCIDATA_27) );
    zdffqb_ PCIDATA_reg_26 ( .CK(PCICLK), .D(PCIDATA_T_26), .Q(PCIDATA_26) );
    zdffqb_ PCIDATA_reg_25 ( .CK(PCICLK), .D(PCIDATA_T_25), .Q(PCIDATA_25) );
    zdffqb_ PCIDATA_reg_24 ( .CK(PCICLK), .D(PCIDATA_T_24), .Q(PCIDATA_24) );
    zdffqb_ PCIDATA_reg_23 ( .CK(PCICLK), .D(PCIDATA_T_23), .Q(PCIDATA_23) );
    zdffqb_ PCIDATA_reg_22 ( .CK(PCICLK), .D(PCIDATA_T_22), .Q(PCIDATA_22) );
    zdffqb_ PCIDATA_reg_21 ( .CK(PCICLK), .D(PCIDATA_T_21), .Q(PCIDATA_21) );
    zdffqb_ PCIDATA_reg_20 ( .CK(PCICLK), .D(PCIDATA_T_20), .Q(PCIDATA_20) );
    zdffqb_ PCIDATA_reg_19 ( .CK(PCICLK), .D(PCIDATA_T_19), .Q(PCIDATA_19) );
    zdffqb_ PCIDATA_reg_18 ( .CK(PCICLK), .D(PCIDATA_T_18), .Q(PCIDATA_18) );
    zdffqb_ PCIDATA_reg_17 ( .CK(PCICLK), .D(PCIDATA_T_17), .Q(PCIDATA_17) );
    zdffqb_ PCIDATA_reg_16 ( .CK(PCICLK), .D(PCIDATA_T_16), .Q(PCIDATA_16) );
    zdffqb_ PCIDATA_reg_15 ( .CK(PCICLK), .D(PCIDATA_T_15), .Q(PCIDATA_15) );
    zdffqb_ PCIDATA_reg_14 ( .CK(PCICLK), .D(PCIDATA_T_14), .Q(PCIDATA_14) );
    zdffqb_ PCIDATA_reg_13 ( .CK(PCICLK), .D(PCIDATA_T_13), .Q(PCIDATA_13) );
    zdffqb_ PCIDATA_reg_12 ( .CK(PCICLK), .D(PCIDATA_T_12), .Q(PCIDATA_12) );
    zdffqb_ PCIDATA_reg_11 ( .CK(PCICLK), .D(PCIDATA_T_11), .Q(PCIDATA_11) );
    zdffqb_ PCIDATA_reg_10 ( .CK(PCICLK), .D(PCIDATA_T_10), .Q(PCIDATA_10) );
    zdffqb_ PCIDATA_reg_9 ( .CK(PCICLK), .D(PCIDATA_T_9), .Q(PCIDATA_9) );
    zdffqb_ PCIDATA_reg_8 ( .CK(PCICLK), .D(PCIDATA_T_8), .Q(PCIDATA_8) );
    zdffqb_ PCIDATA_reg_7 ( .CK(PCICLK), .D(PCIDATA_T_7), .Q(PCIDATA_7) );
    zdffqb_ PCIDATA_reg_6 ( .CK(PCICLK), .D(PCIDATA_T_6), .Q(PCIDATA_6) );
    zdffqb_ PCIDATA_reg_5 ( .CK(PCICLK), .D(PCIDATA_T_5), .Q(PCIDATA_5) );
    zdffqb_ PCIDATA_reg_4 ( .CK(PCICLK), .D(PCIDATA_T_4), .Q(PCIDATA_4) );
    zdffqb_ PCIDATA_reg_3 ( .CK(PCICLK), .D(PCIDATA_T_3), .Q(PCIDATA_3) );
    zdffqb_ PCIDATA_reg_2 ( .CK(PCICLK), .D(PCIDATA_T_2), .Q(PCIDATA_2) );
    zdffqb_ PCIDATA_reg_1 ( .CK(PCICLK), .D(PCIDATA_T_1), .Q(PCIDATA_1) );
    zdffqb_ PCIDATA_reg_0 ( .CK(PCICLK), .D(PCIDATA_T_0), .Q(PCIDATA_0) );
    zdffqrb rptr_reg_8 ( .CK(PCICLK), .D(n_rptr_8), .R(n3024), .Q(rptr_8) );
    zivb U1437 ( .A(rptr_8), .Y(n3104) );
    zdffqrb rptr_reg_7 ( .CK(PCICLK), .D(n_rptr_7), .R(n3029), .Q(rptr_7) );
    zdffqrb rptr_reg_6 ( .CK(PCICLK), .D(n_rptr_6), .R(n3031), .Q(rptr_6) );
    zdffqrb rptr_reg_5 ( .CK(PCICLK), .D(n_rptr_5), .R(n3025), .Q(rptr_5) );
    zdffqrb rptr_reg_4 ( .CK(PCICLK), .D(n_rptr_4), .R(n3025), .Q(rptr_4) );
    zdffqrb rptr_reg_3 ( .CK(PCICLK), .D(n_rptr_3), .R(n3030), .Q(rptr_3) );
    zdffqrb rptr_reg_2 ( .CK(PCICLK), .D(n_rptr_2), .R(n3028), .Q(rptr_2) );
    zdffqrb rptr_reg_0 ( .CK(PCICLK), .D(n_rptr_0), .R(n3026), .Q(rptr_0) );
    zivb U1438 ( .A(rptr_0), .Y(c1328_1) );
    zdffqrb_ RMA_reg_7 ( .CK(PCICLK), .D(rptr_7), .R(n3026), .Q(RMA[7]) );
    zdffqrb_ RMA_reg_5 ( .CK(PCICLK), .D(rptr_5), .R(n3022), .Q(RMA[5]) );
    zdffqrb_ RMA_reg_4 ( .CK(PCICLK), .D(rptr_4), .R(n3023), .Q(RMA[4]) );
    zdffqrb_ RMA_reg_3 ( .CK(PCICLK), .D(rptr_3), .R(n3024), .Q(RMA[3]) );
    zdffqrb_ RMA_reg_0 ( .CK(PCICLK), .D(rptr_0), .R(n3028), .Q(RMA[0]) );
    zdffqrb FSIZE_reg_1 ( .CK(PCICLK), .D(FSIZE1570_1), .R(n3029), .Q(FSIZE_1)
         );
    zivb U1439 ( .A(FSIZE_1), .Y(n3200) );
    zdffqrb FSIZE_reg_0 ( .CK(PCICLK), .D(FSIZE1570_0), .R(n3028), .Q(FSIZE_0)
         );
    zivb U1440 ( .A(FSIZE_0), .Y(n3201) );
    zdffrb RDFF_reg_1 ( .CK(PCICLK), .D(RDFFNXT_1), .R(n3025), .QN(n3068) );
    zdffqrb RDFF_reg_0 ( .CK(PCICLK), .D(RDFFNXT_0), .R(n3029), .Q(RDFFNXT_1)
         );
    zivb U1441 ( .A(RDFFNXT_1), .Y(n3192) );
    zdffqb FFRDPCI_reg_31 ( .CK(PCICLK), .D(FFRDPCI1761_31), .Q(FFRDPCI[31])
         );
    zdffqb FFRDPCI_reg_30 ( .CK(PCICLK), .D(FFRDPCI1761_30), .Q(FFRDPCI[30])
         );
    zdffqb FFRDPCI_reg_29 ( .CK(PCICLK), .D(FFRDPCI1761_29), .Q(FFRDPCI[29])
         );
    zdffqb FFRDPCI_reg_28 ( .CK(PCICLK), .D(FFRDPCI1761_28), .Q(FFRDPCI[28])
         );
    zdffqb FFRDPCI_reg_27 ( .CK(PCICLK), .D(FFRDPCI1761_27), .Q(FFRDPCI[27])
         );
    zdffqb FFRDPCI_reg_26 ( .CK(PCICLK), .D(FFRDPCI1761_26), .Q(FFRDPCI[26])
         );
    zdffqb FFRDPCI_reg_25 ( .CK(PCICLK), .D(FFRDPCI1761_25), .Q(FFRDPCI[25])
         );
    zdffqb FFRDPCI_reg_24 ( .CK(PCICLK), .D(FFRDPCI1761_24), .Q(FFRDPCI[24])
         );
    zdffqb FFRDPCI_reg_23 ( .CK(PCICLK), .D(FFRDPCI1761_23), .Q(FFRDPCI[23])
         );
    zdffqb FFRDPCI_reg_22 ( .CK(PCICLK), .D(FFRDPCI1761_22), .Q(FFRDPCI[22])
         );
    zdffqb FFRDPCI_reg_21 ( .CK(PCICLK), .D(FFRDPCI1761_21), .Q(FFRDPCI[21])
         );
    zdffqb FFRDPCI_reg_20 ( .CK(PCICLK), .D(FFRDPCI1761_20), .Q(FFRDPCI[20])
         );
    zdffqb FFRDPCI_reg_19 ( .CK(PCICLK), .D(FFRDPCI1761_19), .Q(FFRDPCI[19])
         );
    zdffqb FFRDPCI_reg_18 ( .CK(PCICLK), .D(FFRDPCI1761_18), .Q(FFRDPCI[18])
         );
    zdffqb FFRDPCI_reg_17 ( .CK(PCICLK), .D(FFRDPCI1761_17), .Q(FFRDPCI[17])
         );
    zdffqb FFRDPCI_reg_16 ( .CK(PCICLK), .D(FFRDPCI1761_16), .Q(FFRDPCI[16])
         );
    zdffqb FFRDPCI_reg_15 ( .CK(PCICLK), .D(FFRDPCI1761_15), .Q(FFRDPCI[15])
         );
    zdffqb FFRDPCI_reg_14 ( .CK(PCICLK), .D(FFRDPCI1761_14), .Q(FFRDPCI[14])
         );
    zdffqb FFRDPCI_reg_13 ( .CK(PCICLK), .D(FFRDPCI1761_13), .Q(FFRDPCI[13])
         );
    zdffqb FFRDPCI_reg_12 ( .CK(PCICLK), .D(FFRDPCI1761_12), .Q(FFRDPCI[12])
         );
    zdffqb FFRDPCI_reg_11 ( .CK(PCICLK), .D(FFRDPCI1761_11), .Q(FFRDPCI[11])
         );
    zdffqb FFRDPCI_reg_10 ( .CK(PCICLK), .D(FFRDPCI1761_10), .Q(FFRDPCI[10])
         );
    zdffqb FFRDPCI_reg_9 ( .CK(PCICLK), .D(FFRDPCI1761_9), .Q(FFRDPCI[9]) );
    zdffqb FFRDPCI_reg_8 ( .CK(PCICLK), .D(FFRDPCI1761_8), .Q(FFRDPCI[8]) );
    zdffqb FFRDPCI_reg_7 ( .CK(PCICLK), .D(FFRDPCI1761_7), .Q(FFRDPCI[7]) );
    zdffqb FFRDPCI_reg_6 ( .CK(PCICLK), .D(FFRDPCI1761_6), .Q(FFRDPCI[6]) );
    zdffqb FFRDPCI_reg_5 ( .CK(PCICLK), .D(FFRDPCI1761_5), .Q(FFRDPCI[5]) );
    zdffqb FFRDPCI_reg_4 ( .CK(PCICLK), .D(FFRDPCI1761_4), .Q(FFRDPCI[4]) );
    zdffqb FFRDPCI_reg_3 ( .CK(PCICLK), .D(FFRDPCI1761_3), .Q(FFRDPCI[3]) );
    zdffqb FFRDPCI_reg_2 ( .CK(PCICLK), .D(FFRDPCI1761_2), .Q(FFRDPCI[2]) );
    zdffqb FFRDPCI_reg_1 ( .CK(PCICLK), .D(FFRDPCI1761_1), .Q(FFRDPCI[1]) );
    zdffqb FFRDPCI_reg_0 ( .CK(PCICLK), .D(FFRDPCI1761_0), .Q(FFRDPCI[0]) );
    zdffqrb_ TCNT_reg_1 ( .CK(CLK60M), .D(TCNT1958_1), .R(n3025), .Q(n2587) );
    zivb U1442 ( .A(n2587), .Y(n3188) );
    zdffrb ST_BE_reg_1 ( .CK(PCICLK), .D(ST_BE2037_1), .R(n3027), .QN(n3189)
         );
    zdffqrb ST_BE_reg_0 ( .CK(PCICLK), .D(ST_BE2037_0), .R(n3022), .Q(ST_BE_0)
         );
    zivb U1443 ( .A(ST_BE_0), .Y(n3191) );
    zdffqrb END_BE_reg_1 ( .CK(PCICLK), .D(END_BE2076_1), .R(n3029), .Q(
        END_BE_1) );
    zdffqrb END_BE_reg_0 ( .CK(PCICLK), .D(END_BE2076_0), .R(n3027), .Q(
        END_BE_0) );
    zivb U1444 ( .A(END_BE_0), .Y(n3204) );
    zdffqb_ FFRDUSB_reg_31 ( .CK(CLK60M), .D(FFRDUSB2141_31), .Q(FFRDUSB_31)
         );
    zdffqb_ FFRDUSB_reg_30 ( .CK(CLK60M), .D(FFRDUSB2141_30), .Q(FFRDUSB_30)
         );
    zdffqb_ FFRDUSB_reg_29 ( .CK(CLK60M), .D(FFRDUSB2141_29), .Q(FFRDUSB_29)
         );
    zdffqb_ FFRDUSB_reg_28 ( .CK(CLK60M), .D(FFRDUSB2141_28), .Q(FFRDUSB_28)
         );
    zdffqb_ FFRDUSB_reg_27 ( .CK(CLK60M), .D(FFRDUSB2141_27), .Q(FFRDUSB_27)
         );
    zdffqb_ FFRDUSB_reg_26 ( .CK(CLK60M), .D(FFRDUSB2141_26), .Q(FFRDUSB_26)
         );
    zdffqb_ FFRDUSB_reg_25 ( .CK(CLK60M), .D(FFRDUSB2141_25), .Q(FFRDUSB_25)
         );
    zdffqb_ FFRDUSB_reg_24 ( .CK(CLK60M), .D(FFRDUSB2141_24), .Q(FFRDUSB_24)
         );
    zdffqb_ FFRDUSB_reg_23 ( .CK(CLK60M), .D(FFRDUSB2141_23), .Q(FFRDUSB_23)
         );
    zdffqb_ FFRDUSB_reg_22 ( .CK(CLK60M), .D(FFRDUSB2141_22), .Q(FFRDUSB_22)
         );
    zdffqb_ FFRDUSB_reg_21 ( .CK(CLK60M), .D(FFRDUSB2141_21), .Q(FFRDUSB_21)
         );
    zdffqb_ FFRDUSB_reg_20 ( .CK(CLK60M), .D(FFRDUSB2141_20), .Q(FFRDUSB_20)
         );
    zdffqb_ FFRDUSB_reg_19 ( .CK(CLK60M), .D(FFRDUSB2141_19), .Q(FFRDUSB_19)
         );
    zdffqb_ FFRDUSB_reg_18 ( .CK(CLK60M), .D(FFRDUSB2141_18), .Q(FFRDUSB_18)
         );
    zdffqb_ FFRDUSB_reg_17 ( .CK(CLK60M), .D(FFRDUSB2141_17), .Q(FFRDUSB_17)
         );
    zdffqb_ FFRDUSB_reg_16 ( .CK(CLK60M), .D(FFRDUSB2141_16), .Q(FFRDUSB_16)
         );
    zdffqb_ FFRDUSB_reg_15 ( .CK(CLK60M), .D(FFRDUSB2141_15), .Q(FFRDUSB_15)
         );
    zdffqb_ FFRDUSB_reg_14 ( .CK(CLK60M), .D(FFRDUSB2141_14), .Q(FFRDUSB_14)
         );
    zdffqb_ FFRDUSB_reg_13 ( .CK(CLK60M), .D(FFRDUSB2141_13), .Q(FFRDUSB_13)
         );
    zdffqb_ FFRDUSB_reg_12 ( .CK(CLK60M), .D(FFRDUSB2141_12), .Q(FFRDUSB_12)
         );
    zdffqb_ FFRDUSB_reg_11 ( .CK(CLK60M), .D(FFRDUSB2141_11), .Q(FFRDUSB_11)
         );
    zdffqb_ FFRDUSB_reg_10 ( .CK(CLK60M), .D(FFRDUSB2141_10), .Q(FFRDUSB_10)
         );
    zdffqb_ FFRDUSB_reg_9 ( .CK(CLK60M), .D(FFRDUSB2141_9), .Q(FFRDUSB_9) );
    zdffqb_ FFRDUSB_reg_8 ( .CK(CLK60M), .D(FFRDUSB2141_8), .Q(FFRDUSB_8) );
    zdffqb_ FFRDUSB_reg_7 ( .CK(CLK60M), .D(FFRDUSB2141_7), .Q(FFRDUSB_7) );
    zdffqb_ FFRDUSB_reg_6 ( .CK(CLK60M), .D(FFRDUSB2141_6), .Q(FFRDUSB_6) );
    zdffqb_ FFRDUSB_reg_5 ( .CK(CLK60M), .D(FFRDUSB2141_5), .Q(FFRDUSB_5) );
    zdffqb_ FFRDUSB_reg_4 ( .CK(CLK60M), .D(FFRDUSB2141_4), .Q(FFRDUSB_4) );
    zdffqb_ FFRDUSB_reg_3 ( .CK(CLK60M), .D(FFRDUSB2141_3), .Q(FFRDUSB_3) );
    zdffqb_ FFRDUSB_reg_2 ( .CK(CLK60M), .D(FFRDUSB2141_2), .Q(FFRDUSB_2) );
    zdffqb_ FFRDUSB_reg_1 ( .CK(CLK60M), .D(FFRDUSB2141_1), .Q(FFRDUSB_1) );
    zdffqb_ FFRDUSB_reg_0 ( .CK(CLK60M), .D(FFRDUSB2141_0), .Q(FFRDUSB_0) );
    zdffqrb FBE__reg_2 ( .CK(PCICLK), .D(FBE_2296_2), .R(n3031), .Q(FBE_[2])
         );
    zdffqrb FBE__reg_1 ( .CK(PCICLK), .D(FBE_2296_1), .R(n3022), .Q(FBE_[1])
         );
    zdffqrb PROCESS_reg ( .CK(CLK60M), .D(PROCESS2334), .R(n3022), .Q(PROCESS)
         );
    zivb U1445 ( .A(PROCESS), .Y(n3091) );
    zdffqrb PCIWRT_TEST_reg ( .CK(PCICLK), .D(PCIWRT_TEST1184), .R(n3007), .Q(
        PCIWRT_TEST) );
    zdffqrb EOT_2T_reg ( .CK(CLK60M), .D(n3237), .R(n3024), .Q(EOT_2T) );
    zdffqrb_ EOT_PCLK_2T_reg ( .CK(PCICLK), .D(EOT), .R(n3025), .Q(EOT_PCLK_2T
        ) );
    zdffqrb EOT3_2T_reg ( .CK(PCICLK), .D(n3236), .R(n3031), .Q(EOT3_2T) );
    zdffqrb EOT_T_reg ( .CK(CLK60M), .D(EOT_PCLK), .R(n3024), .Q(EOT_T) );
    zdffqrb_ FPOP_T_reg ( .CK(PCICLK), .D(n3235), .R(n3029), .Q(FPOP_T) );
    zdffqrb EOT3_T_reg ( .CK(PCICLK), .D(EOT3_T1447), .R(n3026), .Q(EOT3_T) );
    zivb U1446 ( .A(EOT3_T), .Y(n3205) );
    zdffrb RXPKTEND_T_reg ( .CK(PCICLK), .D(RXPKTEND_T2371), .R(n3022), .QN(
        n3083) );
    zdffqrb_ PIPE_START_T_reg ( .CK(PCICLK), .D(n3234), .R(n3023), .Q(
        PIPE_START_T) );
    zdffqrb_ USBREAD_reg ( .CK(CLK60M), .D(n2952), .R(n3028), .Q(USBREAD) );
    zdffqrb_ RDFF_EQ_WAIT_reg ( .CK(PCICLK), .D(n2949), .R(n3030), .Q(
        RDFF_EQ_WAIT) );
    zdffrb RXPKTEND_reg ( .CK(PCICLK), .D(RXPKTEND2408), .R(n3031), .Q(
        RXPKTEND), .QN(n3082) );
    zdffqrb RXWRT_reg ( .CK(CLK60M), .D(val628_1), .R(n3028), .Q(RXWRT) );
    zdffqrb FPOP_ONCE_reg ( .CK(PCICLK), .D(FPOP_ONCE1612), .R(n3027), .Q(
        FPOP_ONCE) );
    zivb U1447 ( .A(FPOP_ONCE), .Y(n3064) );
    zdffqrb PSH_reg ( .CK(PCICLK), .D(PSH1244), .R(n3030), .Q(PSH) );
    zdffqrb_ PIPE_START_reg ( .CK(PCICLK), .D(PIPE_START1493), .R(n3031), .Q(
        PIPE_START) );
    zdffqrb_ TEST_START_reg ( .CK(PCICLK), .D(TEST_PACKET), .R(n3007), .Q(
        TEST_START) );
    zdffqrb_ LDWPR_2T_reg ( .CK(PCICLK), .D(LDWPR), .R(n3024), .Q(LDWPR_2T) );
    zdffqrb EOT_PCLK_T_reg ( .CK(PCICLK), .D(EOT), .R(n3024), .Q(EOT_PCLK_T)
         );
    znr2b U1448 ( .A(n3068), .B(n3192), .Y(n2949) );
    znr4b U1449 ( .A(n3184), .B(n3185), .C(TESTAD[1]), .D(n3183), .Y(TESTPKTOK
        ) );
    znr2b U1450 ( .A(RXFIFO), .B(n3206), .Y(n2951) );
    znr3b U1451 ( .A(n3187), .B(n3188), .C(n3190), .Y(n2952) );
    znr2b U1452 ( .A(_cell_531_U22_Z_0), .B(n3186), .Y(n2953) );
    znr2b U1453 ( .A(n3199), .B(n3001), .Y(n2954) );
    zaoi21b U1454 ( .A(_cell_531_U22_Z_0), .B(n3066), .C(n3194), .Y(n2955) );
    znr3d U1455 ( .A(n2961), .B(n3085), .C(n3066), .Y(n2956) );
    znr3b U1456 ( .A(FIRSTDW2259), .B(n3189), .C(n3071), .Y(n2957) );
    znr2b U1457 ( .A(n2951), .B(n3000), .Y(n2958) );
    znr2b U1458 ( .A(FIRSTDW2259), .B(n3202), .Y(n2959) );
    znr2b U1459 ( .A(RDFFNXT_1), .B(n3068), .Y(n2960) );
    znr6b U1460 ( .A(rptr_5), .B(rptr_6), .C(rptr_4), .D(rptr_1), .E(rptr_7), 
        .F(n3221), .Y(n2961) );
    znr2b U1461 ( .A(n3113), .B(n3106), .Y(n2962) );
    zoa22b U1462 ( .A(n3109), .B(n3110), .C(n2962), .D(n3108), .Y(n2963) );
    zoa22b U1463 ( .A(n3110), .B(n3112), .C(n2962), .D(n3111), .Y(n2964) );
    znr2b U1464 ( .A(n3075), .B(n3078), .Y(n2965) );
    zoa22b U1465 ( .A(n3115), .B(n3079), .C(n2965), .D(n3114), .Y(n2966) );
    zoa22b U1466 ( .A(n3079), .B(n3117), .C(n2965), .D(n3116), .Y(n2967) );
    zoa22b U1467 ( .A(n3079), .B(n3119), .C(n2965), .D(n3118), .Y(n2968) );
    zoa22b U1468 ( .A(n3079), .B(n3121), .C(n2965), .D(n3120), .Y(n2969) );
    znr2b U1469 ( .A(n3107), .B(n3078), .Y(n2970) );
    zoa22b U1470 ( .A(n3103), .B(n3115), .C(n2970), .D(n3122), .Y(n2971) );
    zoa22b U1471 ( .A(n3103), .B(n3117), .C(n2970), .D(n3123), .Y(n2972) );
    zoa22b U1472 ( .A(n3079), .B(n3125), .C(n2965), .D(n3124), .Y(n2973) );
    zoa22b U1473 ( .A(n3103), .B(n3119), .C(n2970), .D(n3126), .Y(n2974) );
    zoa22b U1474 ( .A(n3103), .B(n3121), .C(n2970), .D(n3127), .Y(n2975) );
    zoa22b U1475 ( .A(n3103), .B(n3125), .C(n2970), .D(n3128), .Y(n2976) );
    zoa22b U1476 ( .A(n3103), .B(n3130), .C(n2970), .D(n3129), .Y(n2977) );
    zoa22b U1477 ( .A(n3103), .B(n3109), .C(n2970), .D(n3131), .Y(n2978) );
    zoa22b U1478 ( .A(n3103), .B(n3112), .C(n2970), .D(n3132), .Y(n2979) );
    znr2b U1479 ( .A(n3077), .B(n3106), .Y(n2980) );
    zoa22b U1480 ( .A(n3115), .B(n3134), .C(n2980), .D(n3133), .Y(n2981) );
    zoa22b U1481 ( .A(n3117), .B(n3134), .C(n2980), .D(n3135), .Y(n2982) );
    zoa22b U1482 ( .A(n3119), .B(n3134), .C(n2980), .D(n3136), .Y(n2983) );
    zoa22b U1483 ( .A(n3121), .B(n3134), .C(n2980), .D(n3137), .Y(n2984) );
    zoa22b U1484 ( .A(n3079), .B(n3130), .C(n2965), .D(n3138), .Y(n2985) );
    zoa22b U1485 ( .A(n3125), .B(n3134), .C(n2980), .D(n3139), .Y(n2986) );
    zoa22b U1486 ( .A(n3130), .B(n3134), .C(n2980), .D(n3140), .Y(n2987) );
    zoa22b U1487 ( .A(n3109), .B(n3134), .C(n2980), .D(n3141), .Y(n2988) );
    zoa22b U1488 ( .A(n3112), .B(n3134), .C(n2980), .D(n3142), .Y(n2989) );
    zoa22b U1489 ( .A(n3110), .B(n3115), .C(n2962), .D(n3143), .Y(n2990) );
    zoa22b U1490 ( .A(n3110), .B(n3117), .C(n2962), .D(n3144), .Y(n2991) );
    zoa22b U1491 ( .A(n3110), .B(n3119), .C(n2962), .D(n3145), .Y(n2992) );
    zoa22b U1492 ( .A(n3110), .B(n3121), .C(n2962), .D(n3146), .Y(n2993) );
    zoa22b U1493 ( .A(n3110), .B(n3125), .C(n2962), .D(n3147), .Y(n2994) );
    zoa22b U1494 ( .A(n3110), .B(n3130), .C(n2962), .D(n3148), .Y(n2995) );
    zoa22b U1495 ( .A(n3109), .B(n3079), .C(n2965), .D(n3149), .Y(n2996) );
    zoa22b U1496 ( .A(n3112), .B(n3079), .C(n2965), .D(n3150), .Y(n2997) );
    znr3b U1497 ( .A(PIPE_START_2T), .B(PIPE_START_T), .C(PIPE_START), .Y(
        n2998) );
    znr3b U1498 ( .A(LDWPR_2T), .B(LDWPR_T), .C(LDWPR), .Y(n2999) );
    znr2b U1499 ( .A(n3100), .B(n3193), .Y(n3000) );
    zaoi211b U1500 ( .A(n3200), .B(n3201), .C(n3074), .D(n3198), .Y(n3001) );
    znr4b U1501 ( .A(FSIZE_0), .B(FSIZE_1), .C(n3096), .D(n3105), .Y(FEMPTY)
         );
    zivb U1502 ( .A(FPUSH), .Y(_cell_531_U22_Z_0) );
    zor2b U1503 ( .A(n3085), .B(n3086), .Y(_cell_531_U41_Z_0) );
    zivb U1504 ( .A(_cell_531_U41_Z_0), .Y(n3199) );
    zdffqrb_ TCNT_reg_0 ( .CK(CLK60M), .D(TCNT1958_0), .R(n3026), .Q(n2586) );
    zivb U1505 ( .A(n2586), .Y(n3190) );
    zdffqrb TESTAD_reg_0 ( .CK(PCICLK), .D(TESTAD1143_0), .R(n3007), .Q(TESTAD
        [0]) );
    zivb U1506 ( .A(TESTAD[0]), .Y(n3183) );
    zdffqrb RCNT_reg_0 ( .CK(CLK60M), .D(RCNT351_0), .R(n3027), .Q(RCNT_0) );
    zivb U1507 ( .A(RCNT_0), .Y(n3102) );
    ziv11b U1508 ( .A(TEST_PACKET), .Y(n3003), .Z(n3004) );
    zivb U1509 ( .A(n3005), .Y(n3232) );
    ziv11b U1510 ( .A(LATCHDAT), .Y(n3005), .Z(n3006) );
    zoa21b U1511 ( .A(ATPG_ENI), .B(n3004), .C(n3027), .Y(n3007) );
    znr3b U1512 ( .A(n3094), .B(n3093), .C(n3098), .Y(FFULL) );
    zaoi21b U1513 ( .A(n3099), .B(n3012), .C(n3041), .Y(n3018) );
    zaoi21b U1514 ( .A(n3099), .B(n3016), .C(n3045), .Y(n3019) );
    zoa21b U1515 ( .A(wptr_6), .B(n3035), .C(n3019), .Y(n3020) );
    ziv11b U1516 ( .A(n3032), .Y(n3021), .Z(n3022) );
    zor2b U1517 ( .A(n3033), .B(ATPG_ENI), .Y(n3032) );
    zivb U1518 ( .A(n3021), .Y(n3024) );
    zivb U1519 ( .A(n3021), .Y(n3023) );
    zdffqrb USBFFTMP_reg_26 ( .CK(CLK60M), .D(USBFFTMP655_26), .R(n3023), .Q(
        USBFFTMP_26) );
    zdffqrb USBFFTMP_reg_15 ( .CK(CLK60M), .D(USBFFTMP655_15), .R(n3029), .Q(
        USBFFTMP_15) );
    zdffqrb END_BE_reg_3 ( .CK(PCICLK), .D(END_BE2076_3), .R(n3022), .Q(
        END_BE_3) );
    zdffqrb USBFFTMP_reg_25 ( .CK(CLK60M), .D(USBFFTMP655_25), .R(n3030), .Q(
        USBFFTMP_25) );
    zdffqrb USBFFTMP_reg_6 ( .CK(CLK60M), .D(USBFFTMP655_6), .R(n3024), .Q(
        USBFFTMP_6) );
    zdffqrb END_BE_reg_2 ( .CK(PCICLK), .D(END_BE2076_2), .R(n3026), .Q(
        END_BE_2) );
    zdffqrb FIRSTDW_reg ( .CK(PCICLK), .D(FIRSTDW2259), .R(n3025), .Q(FIRSTDW)
         );
    zdffrb USBTMP_reg_13 ( .CK(CLK60M), .D(USBTMP396_13), .R(n3030), .QN(n3145
        ) );
    zdffrb USBTMP_reg_16 ( .CK(CLK60M), .D(USBTMP396_16), .R(n3027), .QN(n3142
        ) );
    zdffrb USBTMP_reg_30 ( .CK(CLK60M), .D(USBTMP396_30), .R(n3031), .QN(n3123
        ) );
    zdffrb USBTMP_reg_12 ( .CK(CLK60M), .D(USBTMP396_12), .R(n3023), .QN(n3146
        ) );
    zdffqrb FIFOCNT_reg_0 ( .CK(PCICLK), .D(N_FIFOCNT_0), .R(n3029), .Q(
        FIFOCNT_0) );
    zdffqrb_ WMA_reg_7 ( .CK(PCICLK), .D(wptr_7), .R(n3026), .Q(WMA[7]) );
    zdffqrb_ RMA_reg_8 ( .CK(PCICLK), .D(rptr_8), .R(n3025), .Q(RMA[8]) );
    zdffqrb_ RMA_reg_1 ( .CK(PCICLK), .D(rptr_1), .R(n3028), .Q(RMA[1]) );
    zivb U1520 ( .A(n3021), .Y(n3026) );
    zivb U1521 ( .A(n3021), .Y(n3025) );
    zdffqrb LDWPR_reg ( .CK(PCICLK), .D(LDWPR2000), .R(n3027), .Q(LDWPR) );
    zdffqrb USBFFTMP_reg_10 ( .CK(CLK60M), .D(USBFFTMP655_10), .R(n3022), .Q(
        USBFFTMP_10) );
    zdffqrb USBFFTMP_reg_30 ( .CK(CLK60M), .D(USBFFTMP655_30), .R(n3030), .Q(
        USBFFTMP_30) );
    zdffqrb LDWPR_T_reg ( .CK(PCICLK), .D(LDWPR), .R(n3028), .Q(LDWPR_T) );
    zdffqrb USBFFTMP_reg_14 ( .CK(CLK60M), .D(USBFFTMP655_14), .R(n3024), .Q(
        USBFFTMP_14) );
    zdffqrb USBFFTMP_reg_21 ( .CK(CLK60M), .D(USBFFTMP655_21), .R(n3029), .Q(
        USBFFTMP_21) );
    zdffqrb USBFFTMP_reg_19 ( .CK(CLK60M), .D(USBFFTMP655_19), .R(n3025), .Q(
        USBFFTMP_19) );
    zdffqrb FIFO_OK_reg ( .CK(PCICLK), .D(FIFO_OK1699), .R(n3028), .Q(FIFO_OK)
         );
    zdffrb USBTMP_reg_9 ( .CK(CLK60M), .D(USBTMP396_9), .R(n3029), .QN(n3108)
         );
    zdffrb USBTMP_reg_0 ( .CK(CLK60M), .D(USBTMP396_0), .R(n3023), .QN(n3150)
         );
    zdffrb USBTMP_reg_7 ( .CK(CLK60M), .D(USBTMP396_7), .R(n3027), .QN(n3114)
         );
    zdffrb UPOP_reg ( .CK(CLK60M), .D(USBPOP), .R(n3025), .Q(UPOP), .QN(n3187)
         );
    zdffrb USBTMP_reg_11 ( .CK(CLK60M), .D(USBTMP396_11), .R(n3031), .QN(n3147
        ) );
    zdffrb USBTMP_reg_24 ( .CK(CLK60M), .D(USBTMP396_24), .R(n3031), .QN(n3132
        ) );
    zdffqrb rptr_reg_1 ( .CK(PCICLK), .D(n_rptr_1), .R(n3022), .Q(rptr_1) );
    zdffqrb PIPE_START_2T_reg ( .CK(PCICLK), .D(PIPE_START), .R(n3031), .Q(
        PIPE_START_2T) );
    zdffqrb FBE__reg_3 ( .CK(PCICLK), .D(FBE_2296_3), .R(n3030), .Q(FBE_[3])
         );
    zdffqrb FBE__reg_0 ( .CK(PCICLK), .D(FBE_2296_0), .R(n3026), .Q(FBE_[0])
         );
    zdffqrb_ WMA_reg_8 ( .CK(PCICLK), .D(wptr_8), .R(n3031), .Q(WMA[8]) );
    zdffqrb_ FPUSH_reg ( .CK(PCICLK), .D(FPUSH770), .R(n3027), .Q(FPUSH) );
    zdffqrb_ WMA_reg_5 ( .CK(PCICLK), .D(wptr_5), .R(n3025), .Q(WMA[5]) );
    zdffqrb_ RMA_reg_2 ( .CK(PCICLK), .D(rptr_2), .R(n3023), .Q(RMA[2]) );
    zdffqrb_ RMA_reg_6 ( .CK(PCICLK), .D(rptr_6), .R(n3030), .Q(RMA[6]) );
    zxo2b U1522 ( .A(add_536_carry_8), .B(FIFOCNT_8), .Y(FCOUNT[8]) );
    zan2b U1523 ( .A(FIFOCNT_7), .B(add_536_carry_7), .Y(add_536_carry_8) );
    zxo2b U1524 ( .A(FIFOCNT_7), .B(add_536_carry_7), .Y(FCOUNT[7]) );
    zan2b U1525 ( .A(FIFOCNT_6), .B(add_536_carry_6), .Y(add_536_carry_7) );
    zxo2b U1526 ( .A(FIFOCNT_6), .B(add_536_carry_6), .Y(FCOUNT[6]) );
    zan2b U1527 ( .A(FIFOCNT_5), .B(add_536_carry_5), .Y(add_536_carry_6) );
    zxo2b U1528 ( .A(FIFOCNT_5), .B(add_536_carry_5), .Y(FCOUNT[5]) );
    zan2b U1529 ( .A(FIFOCNT_4), .B(add_536_carry_4), .Y(add_536_carry_5) );
    zxo2b U1530 ( .A(FIFOCNT_4), .B(add_536_carry_4), .Y(FCOUNT[4]) );
    zan2b U1531 ( .A(FIFOCNT_3), .B(add_536_carry_3), .Y(add_536_carry_4) );
    zxo2b U1532 ( .A(FIFOCNT_3), .B(add_536_carry_3), .Y(FCOUNT[3]) );
    zan2b U1533 ( .A(FIFOCNT_2), .B(add_536_carry_2), .Y(add_536_carry_3) );
    zxo2b U1534 ( .A(FIFOCNT_2), .B(add_536_carry_2), .Y(FCOUNT[2]) );
    zan2b U1535 ( .A(FIFOCNT_0), .B(FSIZE_0), .Y(add_536_carry_1) );
    zxo2b U1536 ( .A(FIFOCNT_0), .B(FSIZE_0), .Y(FCOUNT[0]) );
    zinr2b U1537 ( .A(TRST_), .B(BUISTRT), .Y(n3033) );
    zoa21d U1538 ( .A(wptr_7), .B(n3035), .C(n3020), .Y(n3034) );
    zor3b U1539 ( .A(n3010), .B(n3035), .C(n3036), .Y(n3037) );
    zor3b U1540 ( .A(n3012), .B(n3011), .C(n3037), .Y(n3038) );
    zor3b U1541 ( .A(n3014), .B(n3013), .C(n3038), .Y(n3039) );
    zor3b U1542 ( .A(n3016), .B(n3015), .C(n3039), .Y(n3040) );
    zdffrb wptr_reg_8 ( .CK(PCICLK), .D(n3055), .R(n3026), .Q(wptr_8), .QN(
        n3009) );
    zdffrb wptr_reg_7 ( .CK(PCICLK), .D(n3056), .R(n3023), .Q(wptr_7), .QN(
        n3017) );
    zdffrb wptr_reg_6 ( .CK(PCICLK), .D(n3057), .R(n3027), .Q(wptr_6), .QN(
        n3015) );
    zdffrb wptr_reg_5 ( .CK(PCICLK), .D(n3058), .R(n3030), .Q(wptr_5), .QN(
        n3016) );
    zdffrb wptr_reg_4 ( .CK(PCICLK), .D(n3059), .R(n3030), .Q(wptr_4), .QN(
        n3013) );
    zdffrb wptr_reg_3 ( .CK(PCICLK), .D(n3060), .R(n3022), .Q(wptr_3), .QN(
        n3014) );
    zdffrb wptr_reg_2 ( .CK(PCICLK), .D(n3061), .R(n3024), .Q(wptr_2), .QN(
        n3011) );
    zdffrb wptr_reg_1 ( .CK(PCICLK), .D(n3062), .R(n3028), .Q(wptr_1), .QN(
        n3012) );
    zdffrb wptr_reg_0 ( .CK(PCICLK), .D(n3063), .R(n3023), .Q(wptr_0), .QN(
        n3010) );
    zfa1b add_536_U1_1 ( .A(FSIZE_1), .B(FIFOCNT_1), .CI(add_536_carry_1), 
        .CO(add_536_carry_2), .S(FCOUNT[1]) );
    zfa1b r255_U1_0 ( .A(FSIZE_0), .B(_cell_531_U41_Z_0), .CI(n3199), .CO(
        r255_carry_1), .S(FSIZE1554_0) );
    zfa1b r235_U1_5 ( .A(FIFOCNT_5), .B(_cell_531_U22_Z_0), .CI(r235_carry_5), 
        .CO(r235_carry_6), .S(N_FIFOCNT835_5) );
    zfa1b r235_U1_4 ( .A(FIFOCNT_4), .B(_cell_531_U22_Z_0), .CI(r235_carry_4), 
        .CO(r235_carry_5), .S(N_FIFOCNT835_4) );
    zfa1b r235_U1_3 ( .A(FIFOCNT_3), .B(_cell_531_U22_Z_0), .CI(r235_carry_3), 
        .CO(r235_carry_4), .S(N_FIFOCNT835_3) );
    zfa1b r235_U1_2 ( .A(FIFOCNT_2), .B(_cell_531_U22_Z_0), .CI(r235_carry_2), 
        .CO(r235_carry_3), .S(N_FIFOCNT835_2) );
    zfa1b r235_U1_7 ( .A(FIFOCNT_7), .B(_cell_531_U22_Z_0), .CI(r235_carry_7), 
        .CO(r235_carry_8), .S(N_FIFOCNT835_7) );
    zfa1b r235_U1_0 ( .A(FIFOCNT_0), .B(_cell_531_U22_Z_0), .CI(FPUSH), .CO(
        r235_carry_1), .S(N_FIFOCNT835_0) );
    zfa1b r235_U1_6 ( .A(FIFOCNT_6), .B(_cell_531_U22_Z_0), .CI(r235_carry_6), 
        .CO(r235_carry_7), .S(N_FIFOCNT835_6) );
    zfa1b r235_U1_1 ( .A(FIFOCNT_1), .B(_cell_531_U22_Z_0), .CI(r235_carry_1), 
        .CO(r235_carry_2), .S(N_FIFOCNT835_1) );
    zor3b U1543 ( .A(EOT_PCLK_2T), .B(EOT_PCLK_T), .C(EOT), .Y(EOT_PCLK) );
    zoa21d U1544 ( .A(PIPE_START), .B(RDFFNXT_1), .C(n3068), .Y(RDFFNXT_0) );
    zao211b U1545 ( .A(FBE_[0]), .B(n2959), .C(n2957), .D(n3069), .Y(
        FBE_2296_0) );
    zao211b U1546 ( .A(FBE_[1]), .B(n2959), .C(n2957), .D(n3070), .Y(
        FBE_2296_1) );
    zao222b U1547 ( .A(n2957), .B(ST_BE_0), .C(END_BE_2), .D(n3071), .E(FBE_
        [2]), .F(n2959), .Y(FBE_2296_2) );
    zoa21d U1548 ( .A(n3072), .B(n3073), .C(n3074), .Y(PIPE_START1493) );
    zao21d U1549 ( .A(n3232), .B(n3075), .C(n3076), .Y(val628_1) );
    zao222b U1550 ( .A(UCBEO_[1]), .B(n2951), .C(n3000), .D(n3077), .E(n2958), 
        .F(END_BE_1), .Y(END_BE2076_1) );
    zao222b U1551 ( .A(n3000), .B(n3078), .C(UCBEO_[2]), .D(n2951), .E(n2958), 
        .F(END_BE_2), .Y(END_BE2076_2) );
    zao222b U1552 ( .A(n2951), .B(UCBEO_[3]), .C(n3000), .D(n3079), .E(n2958), 
        .F(END_BE_3), .Y(END_BE2076_3) );
    zao222b U1553 ( .A(PCIDATA_0), .B(n3227), .C(TESTDOUT[0]), .D(n3229), .E(
        n3230), .F(USBFFTMP_0), .Y(MDI[0]) );
    zao222b U1554 ( .A(PCIDATA_1), .B(n3080), .C(TESTDOUT[1]), .D(n3229), .E(
        n3081), .F(USBFFTMP_1), .Y(MDI[1]) );
    zao222b U1555 ( .A(PCIDATA_2), .B(n3227), .C(TESTDOUT[2]), .D(n3228), .E(
        n3230), .F(USBFFTMP_2), .Y(MDI[2]) );
    zao222b U1556 ( .A(PCIDATA_3), .B(n3080), .C(TESTDOUT[3]), .D(n3228), .E(
        n3081), .F(USBFFTMP_3), .Y(MDI[3]) );
    zao222b U1557 ( .A(PCIDATA_4), .B(n3227), .C(TESTDOUT[4]), .D(n3228), .E(
        n3230), .F(USBFFTMP_4), .Y(MDI[4]) );
    zao222b U1558 ( .A(PCIDATA_5), .B(n3080), .C(TESTDOUT[5]), .D(n3228), .E(
        n3081), .F(USBFFTMP_5), .Y(MDI[5]) );
    zao222b U1559 ( .A(PCIDATA_6), .B(n3227), .C(TESTDOUT[6]), .D(n3228), .E(
        n3230), .F(USBFFTMP_6), .Y(MDI[6]) );
    zao222b U1560 ( .A(PCIDATA_7), .B(n3080), .C(TESTDOUT[7]), .D(n3228), .E(
        n3081), .F(USBFFTMP_7), .Y(MDI[7]) );
    zao222b U1561 ( .A(PCIDATA_8), .B(n3227), .C(TESTDOUT[8]), .D(n3228), .E(
        n3230), .F(USBFFTMP_8), .Y(MDI[8]) );
    zao222b U1562 ( .A(n3080), .B(PCIDATA_9), .C(n3228), .D(TESTDOUT[9]), .E(
        n3081), .F(USBFFTMP_9), .Y(MDI[9]) );
    zao222b U1563 ( .A(PCIDATA_10), .B(n3080), .C(TESTDOUT[10]), .D(n3228), 
        .E(n3230), .F(USBFFTMP_10), .Y(MDI[10]) );
    zao222b U1564 ( .A(PCIDATA_11), .B(n3227), .C(TESTDOUT[11]), .D(n3228), 
        .E(n3081), .F(USBFFTMP_11), .Y(MDI[11]) );
    zao222b U1565 ( .A(PCIDATA_12), .B(n3080), .C(TESTDOUT[12]), .D(n3228), 
        .E(n3230), .F(USBFFTMP_12), .Y(MDI[12]) );
    zao222b U1566 ( .A(PCIDATA_13), .B(n3227), .C(TESTDOUT[13]), .D(n3229), 
        .E(n3081), .F(USBFFTMP_13), .Y(MDI[13]) );
    zao222b U1567 ( .A(PCIDATA_14), .B(n3080), .C(TESTDOUT[14]), .D(n3229), 
        .E(n3230), .F(USBFFTMP_14), .Y(MDI[14]) );
    zao222b U1568 ( .A(PCIDATA_15), .B(n3227), .C(TESTDOUT[15]), .D(n3229), 
        .E(n3081), .F(USBFFTMP_15), .Y(MDI[15]) );
    zao222b U1569 ( .A(PCIDATA_16), .B(n3080), .C(TESTDOUT[16]), .D(n3229), 
        .E(n3230), .F(USBFFTMP_16), .Y(MDI[16]) );
    zao222b U1570 ( .A(PCIDATA_17), .B(n3227), .C(TESTDOUT[17]), .D(n3229), 
        .E(n3081), .F(USBFFTMP_17), .Y(MDI[17]) );
    zao222b U1571 ( .A(PCIDATA_18), .B(n3080), .C(TESTDOUT[18]), .D(n3004), 
        .E(n3230), .F(USBFFTMP_18), .Y(MDI[18]) );
    zao222b U1572 ( .A(PCIDATA_19), .B(n3227), .C(TESTDOUT[19]), .D(n3004), 
        .E(n3081), .F(USBFFTMP_19), .Y(MDI[19]) );
    zao222b U1573 ( .A(PCIDATA_20), .B(n3080), .C(TESTDOUT[20]), .D(n3004), 
        .E(n3230), .F(USBFFTMP_20), .Y(MDI[20]) );
    zao222b U1574 ( .A(PCIDATA_21), .B(n3227), .C(TESTDOUT[21]), .D(n3004), 
        .E(n3081), .F(USBFFTMP_21), .Y(MDI[21]) );
    zao222b U1575 ( .A(PCIDATA_22), .B(n3080), .C(TESTDOUT[22]), .D(n3004), 
        .E(n3230), .F(USBFFTMP_22), .Y(MDI[22]) );
    zao222b U1576 ( .A(PCIDATA_23), .B(n3227), .C(TESTDOUT[23]), .D(n3004), 
        .E(n3081), .F(USBFFTMP_23), .Y(MDI[23]) );
    zao222b U1577 ( .A(PCIDATA_24), .B(n3080), .C(TESTDOUT[24]), .D(n3004), 
        .E(n3230), .F(USBFFTMP_24), .Y(MDI[24]) );
    zao222b U1578 ( .A(PCIDATA_25), .B(n3227), .C(TESTDOUT[25]), .D(n3229), 
        .E(n3081), .F(USBFFTMP_25), .Y(MDI[25]) );
    zao222b U1579 ( .A(PCIDATA_26), .B(n3080), .C(TESTDOUT[26]), .D(n3004), 
        .E(n3230), .F(USBFFTMP_26), .Y(MDI[26]) );
    zao222b U1580 ( .A(PCIDATA_27), .B(n3227), .C(TESTDOUT[27]), .D(n3229), 
        .E(n3081), .F(USBFFTMP_27), .Y(MDI[27]) );
    zao222b U1581 ( .A(PCIDATA_28), .B(n3080), .C(TESTDOUT[28]), .D(n3004), 
        .E(n3230), .F(USBFFTMP_28), .Y(MDI[28]) );
    zao222b U1582 ( .A(PCIDATA_29), .B(n3227), .C(TESTDOUT[29]), .D(n3229), 
        .E(n3081), .F(USBFFTMP_29), .Y(MDI[29]) );
    zao222b U1583 ( .A(PCIDATA_30), .B(n3080), .C(TESTDOUT[30]), .D(n3004), 
        .E(n3230), .F(USBFFTMP_30), .Y(MDI[30]) );
    zao222b U1584 ( .A(PCIDATA_31), .B(n3227), .C(TESTDOUT[31]), .D(n3229), 
        .E(n3081), .F(USBFFTMP_31), .Y(MDI[31]) );
    zan4b U1585 ( .A(n3089), .B(n3079), .C(PROCESS), .D(RXFIFO), .Y(n3076) );
    zoa21d U1586 ( .A(FPOP_ONCE), .B(n3091), .C(n3000), .Y(n3073) );
    zan4b U1587 ( .A(n3093), .B(n3094), .C(FIFOCNT_1), .D(n3095), .Y(n3092) );
    zor6b U1588 ( .A(FIFOCNT_4), .B(FIFOCNT_2), .C(FIFOCNT_3), .D(FIFOCNT_7), 
        .E(FIFOCNT_5), .F(FIFOCNT_6), .Y(n3097) );
    zor3b U1589 ( .A(FIFOCNT_8), .B(FIFOCNT_0), .C(n3098), .Y(n3105) );
    zind2d U1590 ( .A(TESTPKTOK), .B(TEST_START), .Y(n3186) );
    zao211b U1591 ( .A(FFULL), .B(FPUSH), .C(n3065), .D(n3195), .Y(n3194) );
    zmux21ld U1592 ( .A(n3114), .B(n2966), .S(n3232), .Y(USBTMP396_7) );
    zmux21ld U1593 ( .A(n3127), .B(n2975), .S(n3232), .Y(USBTMP396_28) );
    zmux21ld U1594 ( .A(n3128), .B(n2976), .S(n3232), .Y(USBTMP396_27) );
    zmux21ld U1595 ( .A(n3129), .B(n2977), .S(n3232), .Y(USBTMP396_26) );
    zmux21ld U1596 ( .A(n3131), .B(n2978), .S(n3232), .Y(USBTMP396_25) );
    zmux21ld U1597 ( .A(n3132), .B(n2979), .S(n3232), .Y(USBTMP396_24) );
    zmux21ld U1598 ( .A(n3133), .B(n2981), .S(n3232), .Y(USBTMP396_23) );
    zmux21ld U1599 ( .A(n3135), .B(n2982), .S(n3232), .Y(USBTMP396_22) );
    zmux21ld U1600 ( .A(n3143), .B(n2990), .S(n3232), .Y(USBTMP396_15) );
    zmux21ld U1601 ( .A(n3145), .B(n2992), .S(n3232), .Y(USBTMP396_13) );
    zmux21ld U1602 ( .A(n3147), .B(n2994), .S(n3232), .Y(USBTMP396_11) );
    zmux21ld U1603 ( .A(n3149), .B(n2996), .S(n3232), .Y(USBTMP396_1) );
    zor4b U1604 ( .A(wptr_0), .B(n3009), .C(wptr_1), .D(wptr_7), .Y(n3220) );
    zinr2b U1605 ( .A(EOT_T), .B(EOT_2T), .Y(n3089) );
    zor4b U1606 ( .A(rptr_3), .B(n3104), .C(rptr_0), .D(rptr_2), .Y(n3221) );
    zao211b U1607 ( .A(TDMAEND), .B(n3100), .C(n3092), .D(n3222), .Y(n3072) );
    zor6b U1608 ( .A(wptr_2), .B(wptr_5), .C(wptr_3), .D(wptr_4), .E(wptr_6), 
        .F(n3220), .Y(n3099) );
    zivh U1609 ( .A(val628_1), .Y(n3207) );
    zor3b U1610 ( .A(n2960), .B(RDFF_EQ_WAIT), .C(n2952), .Y(n3223) );
    zmux21ld U1611 ( .A(RCNT_1), .B(RCNT322_1), .S(n3232), .Y(n3213) );
    zmux21ld U1612 ( .A(RCNT_0), .B(n3102), .S(n3006), .Y(n3214) );
    zor3b U1613 ( .A(n3200), .B(n3074), .C(n3198), .Y(n3218) );
    zivh U1614 ( .A(val628_1), .Y(n3233) );
    zbfb U1615 ( .A(PIPE_START), .Y(n3234) );
    zbfb U1616 ( .A(FPOP_T1737), .Y(n3235) );
    zbfb U1617 ( .A(EOT3_T), .Y(n3236) );
    zbfb U1618 ( .A(EOT_T), .Y(n3237) );
endmodule


module TESTDATA ( PCICLK, TEST_PACKET, TESTAD, TESTDOUT );
input  [3:0] TESTAD;
output [31:0] TESTDOUT;
input  PCICLK, TEST_PACKET;
    wire n70, n69, n31, n32, n33, n34, n35, n36, n37, n38, n40, n42, n62, n63, 
        n64, n65, n66, n67, n68;
    zan3b U12 ( .A(TESTAD[0]), .B(TESTAD[1]), .C(n36), .Y(n64) );
    zor2b U13 ( .A(TESTAD[2]), .B(n63), .Y(n65) );
    zivb U14 ( .A(TESTAD[1]), .Y(n63) );
    zivb U15 ( .A(TESTAD[2]), .Y(n68) );
    zor2b U16 ( .A(n32), .B(n69), .Y(TESTDOUT[7]) );
    zivb U17 ( .A(TESTAD[0]), .Y(n66) );
    zivb U18 ( .A(TESTAD[3]), .Y(n67) );
    zor2b U19 ( .A(n64), .B(n37), .Y(n62) );
    zivb U20 ( .A(n40), .Y(TESTDOUT[10]) );
    zivb U21 ( .A(n42), .Y(TESTDOUT[12]) );
    zivb U22 ( .A(n38), .Y(TESTDOUT[13]) );
    zivb U23 ( .A(n40), .Y(TESTDOUT[14]) );
    zivb U24 ( .A(n42), .Y(TESTDOUT[16]) );
    zivb U25 ( .A(n38), .Y(TESTDOUT[17]) );
    zivb U26 ( .A(n38), .Y(TESTDOUT[19]) );
    zivb U27 ( .A(n42), .Y(TESTDOUT[20]) );
    zivb U28 ( .A(n38), .Y(TESTDOUT[21]) );
    zivb U29 ( .A(n38), .Y(TESTDOUT[23]) );
    zivb U30 ( .A(n40), .Y(TESTDOUT[26]) );
    zor2b U31 ( .A(n33), .B(n36), .Y(TESTDOUT[22]) );
    zivb U32 ( .A(n38), .Y(TESTDOUT[31]) );
    znr2b U33 ( .A(TESTAD[3]), .B(n65), .Y(n31) );
    znr3b U34 ( .A(TESTAD[3]), .B(n66), .C(n65), .Y(n32) );
    zaoi211b U35 ( .A(n65), .B(TESTAD[1]), .C(TESTAD[0]), .D(n67), .Y(n33) );
    znr3b U36 ( .A(n67), .B(n66), .C(n65), .Y(n34) );
    znr3b U37 ( .A(TESTAD[1]), .B(n66), .C(n67), .Y(n35) );
    znr2b U38 ( .A(TESTAD[3]), .B(n68), .Y(n36) );
    znr3b U39 ( .A(TESTAD[2]), .B(TESTAD[1]), .C(n67), .Y(n37) );
    ziv11b U40 ( .A(TESTDOUT[9]), .Y(n38), .Z(TESTDOUT[27]) );
    zor2b U41 ( .A(n31), .B(TESTDOUT[7]), .Y(TESTDOUT[9]) );
    ziv11b U42 ( .A(n69), .Y(n40), .Z(TESTDOUT[30]) );
    zor2b U43 ( .A(n33), .B(TESTDOUT[18]), .Y(n69) );
    ziv11b U44 ( .A(n70), .Y(n42), .Z(TESTDOUT[24]) );
    zbfb U45 ( .A(TESTDOUT[5]), .Y(TESTDOUT[3]) );
    zor2b U46 ( .A(n34), .B(TESTDOUT[1]), .Y(TESTDOUT[5]) );
    zbfb U47 ( .A(TESTDOUT[6]), .Y(TESTDOUT[2]) );
    zbfb U48 ( .A(TESTDOUT[8]), .Y(TESTDOUT[0]) );
    zor2b U49 ( .A(n33), .B(n62), .Y(TESTDOUT[8]) );
    zbfb U50 ( .A(TESTDOUT[25]), .Y(TESTDOUT[11]) );
    zor2b U51 ( .A(n31), .B(TESTDOUT[18]), .Y(TESTDOUT[25]) );
    zivb U52 ( .A(n42), .Y(TESTDOUT[28]) );
    zbfb U53 ( .A(TESTDOUT[29]), .Y(TESTDOUT[15]) );
    zor2b U54 ( .A(n31), .B(TESTDOUT[22]), .Y(TESTDOUT[29]) );
    zor3b U55 ( .A(n32), .B(n35), .C(TESTDOUT[22]), .Y(TESTDOUT[1]) );
    zao211b U56 ( .A(n36), .B(TESTAD[0]), .C(n35), .D(n70), .Y(TESTDOUT[6]) );
    zor3b U57 ( .A(n62), .B(n35), .C(n34), .Y(TESTDOUT[4]) );
    zao211b U58 ( .A(n36), .B(TESTAD[1]), .C(n34), .D(TESTDOUT[8]), .Y(n70) );
    zor3b U59 ( .A(n36), .B(n37), .C(n34), .Y(TESTDOUT[18]) );
endmodule


module HS_ACCESS ( SLADDR, SLREAD, RMA, SLAVEMODE, RADDR, DATARDY, FPOP, RD, 
    SLAVE_ACT, FPUSH, WR, PCICLK, TRST_, BIST_RUN, BIST_ERR_S, BIST_RUN_C, 
    FIFO_MDI, MDI, MDO, WMA, WADDR, ASYNCFIFO, BIST_PATTERN, SRAM_WR, SRAM_RUN, 
    SRAM_ADDR, SRAM_SEL, SRAM_RDATA, SRAM_ID, ATPG_CLK, RADDR_ATPG, WADDR_ATPG, 
    MDI_ATPG );
input  [7:0] SLADDR;
input  [8:0] RMA;
input  [31:0] MDO;
input  [8:0] WMA;
output [8:0] WADDR;
input  [31:0] BIST_PATTERN;
input  [1:0] SRAM_ID;
input  [31:0] FIFO_MDI;
input  [8:0] SRAM_ADDR;
output [31:0] MDI_ATPG;
output [31:0] MDI;
output [8:0] RADDR_ATPG;
output [8:0] RADDR;
output [31:0] SRAM_RDATA;
output [8:0] WADDR_ATPG;
input  [1:0] SRAM_SEL;
input  SLREAD, SLAVEMODE, FPOP, SLAVE_ACT, FPUSH, PCICLK, TRST_, BIST_RUN, 
    ASYNCFIFO, SRAM_WR, SRAM_RUN, ATPG_CLK;
output DATARDY, RD, WR, BIST_ERR_S, BIST_RUN_C;
    wire RPOP, BIST_RADDR_6, BIST_WDATA_9, BIST_WDATA734_9, SPAREO6, 
        BIST_WDATA734_21, SRAM_RDATA1309_1, BIST_RDATA_T_8, 
        BIST_RDATA_T1160_21, BIST_RDATA_5, BIST_RDATA1122_9, BIST_RADDR1065_1, 
        BIST_RDATA_13, BISTSM_0, BIST_RDATA_T_31, SRAM_RDATA1309_13, 
        BIST_RDATA_T_16, BIST_WDATA_11, SRAM_RUN_T, BIST_RDATA1122_27, 
        BIST_RDATA1122_12, BIST_WDATA_24, BIST_RDATA_T_23, BIST_RDATA_T1160_6, 
        SRAM_RDATA1309_26, BIST_WDATA_0, BIST_RDATA_26, BISTSMNXT_7, 
        BIST_WDATA734_28, BIST_WADDR677_2, BIST_WDATA734_0, 
        BIST_RDATA_T1160_14, SRAM_W_T, BIST_RDATA1122_0, BIST_WDATA734_14, 
        BIST_RDATA_T_1, BIST_RDATA_T1160_28, SRAM_RDATA1309_8, 
        BIST_RADDRNXT829_2, BIST_WADDRNXT440_7, BIST_RADDR1065_8, BIST_WADDR_3, 
        BIST_WADDR_4, BIST_WDATA_18, BIST_RDATA_T_18, BIST_RDATA1122_29, 
        BIST_RDATA_T_6, BIST_WDATA734_13, BIST_RDATA1122_7, BIST_WADDRNXT440_0, 
        SPAREO0_, BIST_RADDRNXT829_5, BIST_RDATA_21, BIST_WDATA_7, 
        BIST_RDATA_T1160_13, BIST_WDATA734_7, SPAREO8, BIST_WADDR677_5, 
        BIST_RADDR_8, BIST_WDATA_23, BIST_RDATA1122_15, SRAM_RDATA1309_21, 
        BISTSM_7, BIST_RDATA_T1160_1, BIST_RDATA_T_24, BIST_RDATA_T_11, 
        SRAM_RDATA1309_14, BIST_RDATA1122_20, BIST_WDATA_31, BIST_WDATA_16, 
        BIST_RDATA_2, BIST_RDATA_T1160_26, SRAM_RDATA1309_6, BIST_RDATA_14, 
        BIST_RADDR1065_6, BIST_RDATA_28, BIST_WDATA734_26, BIST_RADDR_1, 
        SPAREO1, BIST_WR1405, BIST_RDATA_T1160_8, SRAM_RDATA1309_28, 
        BIST_WDATA_22, BIST_RDATA1122_14, SRAM_RDATA1309_20, 
        BIST_RDATA_T1160_0, BIST_RDATA_T_25, BIST_RDATA_20, BIST_WDATA_6, 
        SPAREO9, BIST_RDATA_T1160_12, BIST_WDATA734_6, BIST_WADDR677_4, 
        SRAM_R_T, BIST_RDATA_T_7, BIST_WDATA734_12, BIST_RD1353, 
        BIST_RDATA1122_6, BIST_WADDRNXT440_1, BIST_RADDRNXT829_4, BIST_WADDR_5, 
        BIST_RDATA_T_19, BIST_RD, BIST_RDATA1122_28, BIST_RADDR_0, 
        WADDR_ATPG1549_0, BIST_RDATA_T1160_9, SRAM_RDATA1309_29, BIST_RDATA_29, 
        BIST_WDATA734_27, SPAREO0, BIST_RDATA_3, BIST_RDATA_T1160_27, 
        SRAM_RDATA1309_7, BIST_WADDRNXT440_8, BIST_RDATA_15, BIST_RADDR1065_7, 
        BISTSM_6, BIST_RDATA_T_10, SRAM_RDATA1309_15, BIST_WDATA_30, 
        BIST_RDATA1122_21, BIST_WDATA_17, BIST_RUNDER, BISTSM_1, 
        BIST_RDATA_T_30, SRAM_RDATA1309_12, BIST_RDATA_T_17, BIST_WDATA_10, 
        BIST_RDATA1122_26, SRAM_RDATA1309_0, BIST_RDATA_T_9, 
        BIST_RDATA_T1160_20, BIST_RDATA_4, BIST_RDATA1122_8, BIST_RADDR1065_0, 
        BIST_RDATA_12, BIST_WDATA_8, SPAREO7, BIST_WDATA734_8, 
        BIST_WDATA734_20, SRAM_W_T1443, BIST_RADDR_7, BIST_WADDR_2, BISTSM_8, 
        BIST_WDATA_19, BIST_RDATA1122_1, BIST_WDATA734_15, BIST_RDATA_T_0, 
        BIST_RDATA_T1160_29, SRAM_RDATA1309_9, BIST_RADDRNXT829_3, 
        BIST_WADDRNXT440_6, BIST_WDATA_1, BIST_RDATA_27, BIST_RFULL, 
        BISTSMNXT_6, BIST_WDATA734_29, BIST_WADDR677_3, BIST_WDATA734_1, 
        BIST_RDATA_T1160_15, BIST_RDATA1122_13, BIST_WDATA_25, BIST_RDATA_T_22, 
        BIST_RDATA_T1160_7, SRAM_RDATA1309_27, BIST_RDATA_T_29, BIST_RADDR_5, 
        BIST_RDATA1122_18, BIST_WFULL, BIST_WDATA734_22, BIST_WADDR677_8, 
        SPAREO5, BIST_RUN_T, BIST_RADDRNXT829_8, BIST_RADDR1065_2, 
        BIST_RDATA_10, BIST_RDATA_6, SRAM_RDATA1309_2, BIST_RDATA_T1160_22, 
        BIST_RDATA1122_24, BIST_WDATA_12, BISTSM_3, BIST_RDATA_T_15, 
        SRAM_RDATA1309_10, SRAM_RDATA1309_25, BIST_RDATA_T_20, 
        BIST_RDATA_T1160_5, BIST_WDATA_27, BIST_RDATA1122_11, BIST_WDATA734_3, 
        BIST_RDATA_T1160_17, BIST_REMPTY, BISTSMNXT_4, BIST_WADDR677_1, 
        BIST_RDATA_T1160_30, BIST_RDATA_25, BIST_RD_T1359, BIST_WDATA_3, 
        BIST_RDATA_19, BIST_WADDRNXT440_4, BIST_RUN_C346, BIST_RADDRNXT829_1, 
        BIST_RDATA_T_2, BIST_WDATA734_30, BIST_RDATA1122_3, BIST_WDATA734_17, 
        BIST_WADDR_0, SRAM_RDATA1309_19, SRAM_R_T1481, BIST_WADDR_7, 
        BIST_RADDRNXT829_6, BIST_WADDRNXT440_3, BIST_WDATA734_10, BIST_RDATA_8, 
        BIST_RDATA1122_4, BIST_RDATA_T_5, BIST_WADDR677_6, BISTSMNXT_3, 
        BIST_WDATA734_4, BIST_RDATA_T1160_10, BIST_WDATA_4, BIST_RDATA_22, 
        BIST_RDATA_T1160_2, BIST_RDATA_T_27, SRAM_RDATA1309_22, 
        BIST_RDATA1122_16, BIST_RDATA1122_31, BIST_WDATA_20, BIST_WDATA_15, 
        BIST_RDATA1122_23, BISTSM_4, SRAM_RDATA1309_17, BIST_RDATA_T_12, 
        SRAM_RDATA1309_30, BIST_RDATA_17, BIST_RADDR1065_5, BIST_RDATA_30, 
        BIST_RDATA_T1160_25, SRAM_RDATA1309_5, BIST_WDATA734_19, BIST_RDATA_1, 
        SPAREO2, BIST_RDATA_T1160_19, BIST_WDATA734_25, BIST_WR, BIST_WDATA_29, 
        BIST_RADDR_2, BIST_RDATA_T1160_3, BIST_RDATA_T_26, SRAM_RDATA1309_23, 
        BIST_RDATA1122_17, BIST_CMP, BIST_RDATA1122_30, BIST_WDATA_21, 
        BIST_WADDR677_7, BISTSMNXT_2, BIST_WDATA734_5, BIST_RDATA_T1160_11, 
        BIST_WUNDER, BIST_WDATA_5, BIST_RDATA_23, BIST_RADDRNXT829_7, 
        BIST_WADDRNXT440_2, BIST_WDATA734_11, BIST_RDATA_9, BIST_RDATA1122_5, 
        BIST_RDATA_T_4, BIST_ERR_S1235, BIST_WADDR_6, BIST_WDATA_28, 
        BIST_RADDR_3, BIST_RDATA_T1160_18, SPAREO3, BIST_WDATA734_24, SPAREO1_, 
        BIST_RDATA_16, BIST_RADDR1065_4, BIST_RDATA_31, BIST_RDATA_T1160_24, 
        SRAM_RDATA1309_4, BIST_WDATA734_18, BIST_RDATA_0, BIST_WDATA_14, 
        BIST_RDATA1122_22, BISTSM_5, SRAM_RDATA1309_16, RPOP187, 
        BIST_RDATA_T_13, SRAM_RDATA1309_31, BIST_RDATA1122_25, BIST_WADDR_8, 
        BIST_WDATA_13, BISTSM_2, BIST_RDATA_T_14, SRAM_RDATA1309_11, 
        BIST_RADDR1065_3, BIST_RDATA_11, BIST_RDATA_7, SRAM_RDATA1309_3, 
        BIST_RDATA_T1160_23, BIST_WDATA734_23, SPAREO4, BIST_RDATA_T_28, 
        BIST_RADDR_4, BIST_RDATA1122_19, BIST_RD_T, BIST_WADDR_1, 
        SRAM_RDATA1309_18, BIST_WADDRNXT440_5, BIST_RDATA_18, 
        BIST_RADDRNXT829_0, BIST_WDATA734_31, BIST_RDATA_T_3, BIST_RDATA1122_2, 
        BIST_WDATA734_16, BIST_RDATA_T1160_16, BIST_WDATA734_2, BISTSMNXT_5, 
        BIST_RDATA_T1160_31, BIST_WADDR677_0, BIST_RDATA_24, BIST_WDATA_2, 
        SRAM_RDATA1309_24, BIST_RDATA_T_21, BIST_RDATA_T1160_4, BIST_WDATA_26, 
        BIST_RDATA1122_10, n1736, n1740, n1950, n1951, n1952, n1953, n1954, 
        n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, 
        n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, 
        n1975, n1976, n1977, n1978, n1979, n1980, r133_carry_8, r133_carry_1, 
        r133_carry_7, r133_carry_6, r133_carry_2, r133_carry_5, r133_carry_4, 
        r133_carry_3, r143_carry_8, r143_carry_1, r143_carry_7, r143_carry_6, 
        r143_carry_2, r143_carry_5, r143_carry_4, r143_carry_3, n1981, n1982, 
        n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
        n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
        n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
        n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
        n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
        n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
        n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
        n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
        n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
        n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
        n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
        n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
        n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
        n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
        n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
        n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
        n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
        n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
        n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
        n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
        n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
        n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
        n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
        n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, 
        n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, 
        n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, 
        n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, 
        n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
        n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
        n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
        n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, 
        n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, 
        n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, 
        n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, 
        n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, 
        n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, 
        n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, 
        n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, 
        n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, 
        n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, 
        n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, 
        n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
        n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, 
        n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, 
        n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, 
        n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, 
        n2443, n2444, _cell_830_U14_Z_0, _cell_830_U3_Z_0, n2445, n2446;
    zoai21b SPARE685 ( .A(SPAREO1), .B(n1958), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE682 ( .A(SPAREO0), .B(BIST_RFULL), .C(SPAREO1_), .D(1'b0), 
        .Y(SPAREO2) );
    zaoi211b SPARE683 ( .A(SPAREO4), .B(BIST_WFULL), .C(SPAREO6), .D(
        BIST_REMPTY), .Y(SPAREO8) );
    zoai21b SPARE684 ( .A(SPAREO0), .B(SPAREO8), .C(BIST_WUNDER), .Y(SPAREO9)
         );
    znr3b SPARE686 ( .A(SPAREO2), .B(BIST_RUNDER), .C(SPAREO0_), .Y(SPAREO4)
         );
    zivb SPARE688 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE681 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    znd3b SPARE689 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE680 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE687 ( .A(SPAREO4), .Y(SPAREO5) );
    zoai21b U651 ( .A(n2271), .B(n2233), .C(n2382), .Y(n2298) );
    zor2b U652 ( .A(BISTSMNXT_2), .B(BISTSM_0), .Y(n2233) );
    zao21b U653 ( .A(BIST_RFULL), .B(n2258), .C(n2214), .Y(n2257) );
    zivb U654 ( .A(n2257), .Y(n2382) );
    zan3b U655 ( .A(BISTSM_7), .B(n2206), .C(n2268), .Y(n2208) );
    zan2b U656 ( .A(BIST_RFULL), .B(n2187), .Y(n2186) );
    zxo3b r133_U1_8 ( .A(BIST_WADDR_8), .B(_cell_830_U14_Z_0), .C(r133_carry_8
        ), .Y(BIST_WADDRNXT440_8) );
    zoai21b U657 ( .A(n2238), .B(BIST_WUNDER), .C(_cell_830_U14_Z_0), .Y(n2193
        ) );
    zor2b U658 ( .A(n2190), .B(n2235), .Y(n2192) );
    zxo3b r143_U1_8 ( .A(BIST_RADDR_8), .B(_cell_830_U3_Z_0), .C(r143_carry_8), 
        .Y(BIST_RADDRNXT829_8) );
    zor2b U659 ( .A(n2256), .B(n1960), .Y(n2201) );
    zor2b U660 ( .A(n1960), .B(n2256), .Y(n2199) );
    znd8b U661 ( .A(n2309), .B(n2310), .C(n2311), .D(n2312), .E(n2313), .F(
        n2314), .G(n2315), .H(n2316), .Y(n2308) );
    zxo2b U662 ( .A(n2343), .B(BIST_RDATA_T_16), .Y(n2309) );
    zivb U663 ( .A(MDO[16]), .Y(n2343) );
    zxo2b U664 ( .A(n2344), .B(BIST_RDATA_T_22), .Y(n2310) );
    zivb U665 ( .A(MDO[22]), .Y(n2344) );
    zxo2b U666 ( .A(n2345), .B(BIST_RDATA_T_3), .Y(n2311) );
    zivb U667 ( .A(MDO[3]), .Y(n2345) );
    zxo2b U668 ( .A(n2346), .B(BIST_RDATA_T_8), .Y(n2312) );
    zivb U669 ( .A(MDO[8]), .Y(n2346) );
    zxo2b U670 ( .A(n2347), .B(BIST_RDATA_T_30), .Y(n2313) );
    zivb U671 ( .A(MDO[30]), .Y(n2347) );
    zxo2b U672 ( .A(n2348), .B(BIST_RDATA_T_15), .Y(n2314) );
    zivb U673 ( .A(MDO[15]), .Y(n2348) );
    zxo2b U674 ( .A(n2349), .B(BIST_RDATA_T_10), .Y(n2315) );
    zivb U675 ( .A(MDO[10]), .Y(n2349) );
    zxo2b U676 ( .A(n2350), .B(BIST_RDATA_T_28), .Y(n2316) );
    zivb U677 ( .A(MDO[28]), .Y(n2350) );
    znd8b U678 ( .A(n2300), .B(n2301), .C(n2302), .D(n2303), .E(n2304), .F(
        n2305), .G(n2306), .H(n2307), .Y(n2299) );
    zxo2b U679 ( .A(n2335), .B(BIST_RDATA_T_9), .Y(n2300) );
    zivb U680 ( .A(MDO[9]), .Y(n2335) );
    zxo2b U681 ( .A(n2336), .B(BIST_RDATA_T_1), .Y(n2301) );
    zivb U682 ( .A(MDO[1]), .Y(n2336) );
    zxo2b U683 ( .A(n2337), .B(BIST_RDATA_T_24), .Y(n2302) );
    zivb U684 ( .A(MDO[24]), .Y(n2337) );
    zxo2b U685 ( .A(n2338), .B(BIST_RDATA_T_27), .Y(n2303) );
    zivb U686 ( .A(MDO[27]), .Y(n2338) );
    zxo2b U687 ( .A(n2339), .B(BIST_RDATA_T_7), .Y(n2304) );
    zivb U688 ( .A(MDO[7]), .Y(n2339) );
    zxo2b U689 ( .A(n2340), .B(BIST_RDATA_T_21), .Y(n2305) );
    zivb U690 ( .A(MDO[21]), .Y(n2340) );
    zxo2b U691 ( .A(n2341), .B(BIST_RDATA_T_4), .Y(n2306) );
    zivb U692 ( .A(MDO[4]), .Y(n2341) );
    zxo2b U693 ( .A(n2342), .B(BIST_RDATA_T_29), .Y(n2307) );
    zivb U694 ( .A(MDO[29]), .Y(n2342) );
    znd8b U695 ( .A(n2327), .B(n2328), .C(n2329), .D(n2330), .E(n2331), .F(
        n2332), .G(n2333), .H(n2334), .Y(n2326) );
    zxo2b U696 ( .A(n2359), .B(BIST_RDATA_T_13), .Y(n2327) );
    zivb U697 ( .A(MDO[13]), .Y(n2359) );
    zxo2b U698 ( .A(n2360), .B(BIST_RDATA_T_6), .Y(n2328) );
    zivb U699 ( .A(MDO[6]), .Y(n2360) );
    zxo2b U700 ( .A(n2361), .B(BIST_RDATA_T_19), .Y(n2329) );
    zivb U701 ( .A(MDO[19]), .Y(n2361) );
    zxo2b U702 ( .A(n2362), .B(BIST_RDATA_T_14), .Y(n2330) );
    zivb U703 ( .A(MDO[14]), .Y(n2362) );
    zxo2b U704 ( .A(n2363), .B(BIST_RDATA_T_31), .Y(n2331) );
    zivb U705 ( .A(MDO[31]), .Y(n2363) );
    zxo2b U706 ( .A(n2364), .B(BIST_RDATA_T_11), .Y(n2332) );
    zivb U707 ( .A(MDO[11]), .Y(n2364) );
    zxo2b U708 ( .A(n2365), .B(BIST_RDATA_T_17), .Y(n2333) );
    zivb U709 ( .A(MDO[17]), .Y(n2365) );
    zxo2b U710 ( .A(n2366), .B(BIST_RDATA_T_26), .Y(n2334) );
    zivb U711 ( .A(MDO[26]), .Y(n2366) );
    znd8b U712 ( .A(n2318), .B(n2319), .C(n2320), .D(n2321), .E(n2322), .F(
        n2323), .G(n2324), .H(n2325), .Y(n2317) );
    zxo2b U713 ( .A(n2351), .B(BIST_RDATA_T_2), .Y(n2318) );
    zivb U714 ( .A(MDO[2]), .Y(n2351) );
    zxo2b U715 ( .A(n2352), .B(BIST_RDATA_T_23), .Y(n2319) );
    zivb U716 ( .A(MDO[23]), .Y(n2352) );
    zxo2b U717 ( .A(n2353), .B(BIST_RDATA_T_18), .Y(n2320) );
    zivb U718 ( .A(MDO[18]), .Y(n2353) );
    zxo2b U719 ( .A(n2354), .B(BIST_RDATA_T_12), .Y(n2321) );
    zivb U720 ( .A(MDO[12]), .Y(n2354) );
    zxo2b U721 ( .A(n2355), .B(BIST_RDATA_T_25), .Y(n2322) );
    zivb U722 ( .A(MDO[25]), .Y(n2355) );
    zxo2b U723 ( .A(n2356), .B(BIST_RDATA_T_0), .Y(n2323) );
    zivb U724 ( .A(MDO[0]), .Y(n2356) );
    zxo2b U725 ( .A(n2357), .B(BIST_RDATA_T_5), .Y(n2324) );
    zivb U726 ( .A(MDO[5]), .Y(n2357) );
    zxo2b U727 ( .A(n2358), .B(BIST_RDATA_T_20), .Y(n2325) );
    zivb U728 ( .A(MDO[20]), .Y(n2358) );
    zmux21lb U729 ( .A(n2207), .B(n2205), .S(BISTSM_7), .Y(n2248) );
    zan2b U730 ( .A(BISTSM_8), .B(n1972), .Y(n2207) );
    zan2b U731 ( .A(BIST_REMPTY), .B(n2206), .Y(n2205) );
    zivb U732 ( .A(n2231), .Y(n2268) );
    zmux21lb U733 ( .A(n2290), .B(n2291), .S(n1961), .Y(n2261) );
    zmux21lb U734 ( .A(n2277), .B(n2278), .S(n2281), .Y(n2245) );
    zor2b U735 ( .A(BISTSM_5), .B(n2016), .Y(n2224) );
    zmux21lb U736 ( .A(n2290), .B(n2291), .S(n2292), .Y(n2262) );
    zmux21lb U737 ( .A(n2277), .B(n2278), .S(n2280), .Y(n2244) );
    zmux21lb U738 ( .A(n2290), .B(n2291), .S(n2294), .Y(n2264) );
    zan2b U739 ( .A(BISTSM_7), .B(BIST_WUNDER), .Y(n2198) );
    zmux21lb U740 ( .A(n2266), .B(n2267), .S(BIST_WADDR_8), .Y(n2255) );
    zor2b U741 ( .A(n2182), .B(n2162), .Y(n2266) );
    zor2b U742 ( .A(BIST_WADDR_7), .B(ASYNCFIFO), .Y(n2267) );
    zmux21lb U743 ( .A(n2204), .B(n2202), .S(BIST_RADDR_8), .Y(n2229) );
    zan2b U744 ( .A(BIST_RADDR_7), .B(ASYNCFIFO), .Y(n2204) );
    zan2b U745 ( .A(n2162), .B(n2203), .Y(n2202) );
    zmux21lb U746 ( .A(n2277), .B(n2278), .S(n2282), .Y(n2246) );
    zor2b U747 ( .A(n2020), .B(n2259), .Y(n2374) );
    zmux21lb U748 ( .A(n2290), .B(n2291), .S(n2293), .Y(n2263) );
    zor2b U749 ( .A(n2240), .B(n2020), .Y(n2370) );
    zmux21lb U750 ( .A(n2277), .B(n2278), .S(n2279), .Y(n2243) );
    zor2b U751 ( .A(BISTSMNXT_5), .B(BISTSMNXT_7), .Y(n2273) );
    zoai21b U752 ( .A(BISTSMNXT_4), .B(n2233), .C(n2236), .Y(n2371) );
    zivb U753 ( .A(n2371), .Y(n2237) );
    zoai21b U754 ( .A(BIST_WFULL), .B(n2234), .C(n2241), .Y(n2240) );
    zor2b U755 ( .A(BIST_WUNDER), .B(n2187), .Y(n2241) );
    zivb U756 ( .A(n2241), .Y(n2367) );
    zor2b U757 ( .A(n2178), .B(n2278), .Y(n2291) );
    zor2b U758 ( .A(n2368), .B(n2022), .Y(n2290) );
    zoa22b U759 ( .A(BIST_REMPTY), .B(n2195), .C(BIST_RFULL), .D(n2196), .Y(
        n2194) );
    zor2b U760 ( .A(BIST_REMPTY), .B(n2187), .Y(n2258) );
    zor2b U761 ( .A(BIST_RFULL), .B(n2214), .Y(n2022) );
    zivb U762 ( .A(n2022), .Y(n2284) );
    zmux21lb U763 ( .A(n1956), .B(n1955), .S(BIST_RFULL), .Y(n2196) );
    zor2b U764 ( .A(BISTSMNXT_6), .B(BISTSMNXT_7), .Y(n2191) );
    zivb U765 ( .A(n2190), .Y(n2238) );
    zor2b U766 ( .A(BISTSMNXT_4), .B(BISTSMNXT_2), .Y(n2189) );
    zxo2b U767 ( .A(SRAM_SEL[1]), .B(SRAM_ID[1]), .Y(n2211) );
    zxo2b U768 ( .A(SRAM_SEL[0]), .B(SRAM_ID[0]), .Y(n2212) );
    zivb U769 ( .A(n2195), .Y(BISTSMNXT_7) );
    zmux21lb U770 ( .A(n2208), .B(n1957), .S(BIST_REMPTY), .Y(n2195) );
    zao22b U771 ( .A(BIST_RFULL), .B(n1956), .C(n1957), .D(n2011), .Y(
        BISTSMNXT_6) );
    zao22b U772 ( .A(n1954), .B(BIST_REMPTY), .C(n1955), .D(n2009), .Y(
        BISTSMNXT_4) );
    zao22b U773 ( .A(n1953), .B(BIST_RFULL), .C(n1954), .D(n2011), .Y(
        BISTSMNXT_3) );
    zivb U774 ( .A(BISTSMNXT_3), .Y(n2278) );
    zao22b U775 ( .A(n1953), .B(n2009), .C(n2010), .D(BIST_REMPTY), .Y(
        BISTSMNXT_2) );
    zivb U776 ( .A(n2011), .Y(BIST_REMPTY) );
    zivb U777 ( .A(BISTSMNXT_2), .Y(n2368) );
    zor2b U778 ( .A(BISTSM_7), .B(BISTSM_8), .Y(n2223) );
    zmux21lb U779 ( .A(n2271), .B(n2186), .S(BISTSM_0), .Y(n2270) );
    zivb U780 ( .A(n2258), .Y(n2271) );
    zivb U781 ( .A(n2223), .Y(n2295) );
    zor2b U782 ( .A(BISTSM_1), .B(n2223), .Y(n2225) );
    zmux21lb U783 ( .A(n1972), .B(n2009), .S(BISTSM_0), .Y(n2269) );
    zivb U784 ( .A(n2230), .Y(n2296) );
    zcx2b U785 ( .A(n2181), .B(n2193), .C(BIST_WADDRNXT440_8), .D(n2192), .Y(
        n2170) );
    zan2b U786 ( .A(n2163), .B(n2171), .Y(BIST_WADDR677_6) );
    zao22b U787 ( .A(n2376), .B(BIST_WADDR_6), .C(BIST_WADDRNXT440_6), .D(
        n2192), .Y(n2171) );
    zivb U788 ( .A(n2171), .Y(n2280) );
    zan2b U789 ( .A(n2163), .B(n2172), .Y(BIST_WADDR677_5) );
    zao22b U790 ( .A(n2376), .B(BIST_WADDR_5), .C(BIST_WADDRNXT440_5), .D(
        n2192), .Y(n2172) );
    zan2b U791 ( .A(n2163), .B(n2173), .Y(BIST_WADDR677_4) );
    zao22b U792 ( .A(n2376), .B(BIST_WADDR_4), .C(BIST_WADDRNXT440_4), .D(
        n2192), .Y(n2173) );
    zivb U793 ( .A(n2173), .Y(n2281) );
    zan2b U794 ( .A(n2163), .B(n2174), .Y(BIST_WADDR677_3) );
    zao22b U795 ( .A(n2376), .B(BIST_WADDR_3), .C(BIST_WADDRNXT440_3), .D(
        n2192), .Y(n2174) );
    zan2b U796 ( .A(n2163), .B(n2175), .Y(BIST_WADDR677_2) );
    zao22b U797 ( .A(n2376), .B(BIST_WADDR_2), .C(BIST_WADDRNXT440_2), .D(
        n2192), .Y(n2175) );
    zivb U798 ( .A(n2175), .Y(n2282) );
    zan2b U799 ( .A(n2163), .B(n2176), .Y(BIST_WADDR677_1) );
    zao22b U800 ( .A(n2376), .B(BIST_WADDR_1), .C(BIST_WADDRNXT440_1), .D(
        n2192), .Y(n2176) );
    zan2b U801 ( .A(n2163), .B(n2177), .Y(BIST_WADDR677_0) );
    zao22b U802 ( .A(n2376), .B(BIST_WADDR_0), .C(BIST_WADDRNXT440_0), .D(
        n2192), .Y(n2177) );
    zivb U803 ( .A(n2193), .Y(n2376) );
    zivb U804 ( .A(n2177), .Y(n2279) );
    zcx2b U805 ( .A(n2200), .B(n2201), .C(BIST_RADDRNXT829_8), .D(n2199), .Y(
        n2160) );
    zivb U806 ( .A(ASYNCFIFO), .Y(n2162) );
    zan2b U807 ( .A(n2163), .B(n2164), .Y(BIST_RADDR1065_6) );
    zao22b U808 ( .A(n2375), .B(BIST_RADDR_6), .C(BIST_RADDRNXT829_6), .D(
        n2199), .Y(n2164) );
    zivb U809 ( .A(n2164), .Y(n2292) );
    zan2b U810 ( .A(n2163), .B(n2165), .Y(BIST_RADDR1065_5) );
    zao22b U811 ( .A(n2375), .B(BIST_RADDR_5), .C(BIST_RADDRNXT829_5), .D(
        n2199), .Y(n2165) );
    zan2b U812 ( .A(n2163), .B(n2166), .Y(BIST_RADDR1065_4) );
    zao22b U813 ( .A(n2375), .B(BIST_RADDR_4), .C(BIST_RADDRNXT829_4), .D(
        n2199), .Y(n2166) );
    zivb U814 ( .A(n2166), .Y(n2293) );
    zan2b U815 ( .A(n2163), .B(n2167), .Y(BIST_RADDR1065_3) );
    zao22b U816 ( .A(n2375), .B(BIST_RADDR_3), .C(BIST_RADDRNXT829_3), .D(
        n2199), .Y(n2167) );
    zan2b U817 ( .A(n2163), .B(n2168), .Y(BIST_RADDR1065_2) );
    zao22b U818 ( .A(n2375), .B(BIST_RADDR_2), .C(BIST_RADDRNXT829_2), .D(
        n2199), .Y(n2168) );
    zivb U819 ( .A(n2168), .Y(n2294) );
    zan2b U820 ( .A(n2163), .B(n2169), .Y(BIST_RADDR1065_1) );
    zao22b U821 ( .A(n2375), .B(BIST_RADDR_1), .C(BIST_RADDRNXT829_1), .D(
        n2199), .Y(n2169) );
    zoai21b U822 ( .A(n1961), .B(n2161), .C(n2159), .Y(BIST_RADDR1065_0) );
    zivb U823 ( .A(n2201), .Y(n2375) );
    zivb U824 ( .A(n2159), .Y(n2247) );
    zor2b U825 ( .A(BISTSM_7), .B(n2195), .Y(n2159) );
    zivb U826 ( .A(n2161), .Y(n2163) );
    zmux21hb U827 ( .A(SRAM_RDATA[31]), .B(MDO[31]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_31) );
    zmux21hb U828 ( .A(SRAM_RDATA[30]), .B(MDO[30]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_30) );
    zmux21hb U829 ( .A(SRAM_RDATA[29]), .B(MDO[29]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_29) );
    zmux21hb U830 ( .A(SRAM_RDATA[28]), .B(MDO[28]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_28) );
    zmux21hb U831 ( .A(SRAM_RDATA[27]), .B(MDO[27]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_27) );
    zmux21hb U832 ( .A(SRAM_RDATA[26]), .B(MDO[26]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_26) );
    zmux21hb U833 ( .A(SRAM_RDATA[25]), .B(MDO[25]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_25) );
    zmux21hb U834 ( .A(SRAM_RDATA[24]), .B(MDO[24]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_24) );
    zmux21hb U835 ( .A(SRAM_RDATA[23]), .B(MDO[23]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_23) );
    zmux21hb U836 ( .A(SRAM_RDATA[22]), .B(MDO[22]), .S(n1980), .Y(
        SRAM_RDATA1309_22) );
    zmux21hb U837 ( .A(SRAM_RDATA[21]), .B(MDO[21]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_21) );
    zmux21hb U838 ( .A(SRAM_RDATA[20]), .B(MDO[20]), .S(n1980), .Y(
        SRAM_RDATA1309_20) );
    zmux21hb U839 ( .A(SRAM_RDATA[19]), .B(MDO[19]), .S(n1980), .Y(
        SRAM_RDATA1309_19) );
    zmux21hb U840 ( .A(SRAM_RDATA[18]), .B(MDO[18]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_18) );
    zmux21hb U841 ( .A(SRAM_RDATA[17]), .B(MDO[17]), .S(n1980), .Y(
        SRAM_RDATA1309_17) );
    zmux21hb U842 ( .A(SRAM_RDATA[16]), .B(MDO[16]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_16) );
    zmux21hb U843 ( .A(SRAM_RDATA[15]), .B(MDO[15]), .S(n1980), .Y(
        SRAM_RDATA1309_15) );
    zmux21hb U844 ( .A(SRAM_RDATA[14]), .B(MDO[14]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_14) );
    zmux21hb U845 ( .A(SRAM_RDATA[13]), .B(MDO[13]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_13) );
    zmux21hb U846 ( .A(SRAM_RDATA[12]), .B(MDO[12]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_12) );
    zmux21hb U847 ( .A(SRAM_RDATA[11]), .B(MDO[11]), .S(n1980), .Y(
        SRAM_RDATA1309_11) );
    zmux21hb U848 ( .A(SRAM_RDATA[10]), .B(MDO[10]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_10) );
    zmux21hb U849 ( .A(SRAM_RDATA[9]), .B(MDO[9]), .S(n1980), .Y(
        SRAM_RDATA1309_9) );
    zmux21hb U850 ( .A(SRAM_RDATA[8]), .B(MDO[8]), .S(n1980), .Y(
        SRAM_RDATA1309_8) );
    zmux21hb U851 ( .A(SRAM_RDATA[7]), .B(MDO[7]), .S(n1980), .Y(
        SRAM_RDATA1309_7) );
    zmux21hb U852 ( .A(SRAM_RDATA[6]), .B(MDO[6]), .S(n1980), .Y(
        SRAM_RDATA1309_6) );
    zmux21hb U853 ( .A(SRAM_RDATA[5]), .B(MDO[5]), .S(n1980), .Y(
        SRAM_RDATA1309_5) );
    zmux21hb U854 ( .A(SRAM_RDATA[4]), .B(MDO[4]), .S(n1980), .Y(
        SRAM_RDATA1309_4) );
    zmux21hb U855 ( .A(SRAM_RDATA[3]), .B(MDO[3]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_3) );
    zmux21hb U856 ( .A(SRAM_RDATA[2]), .B(MDO[2]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_2) );
    zmux21hb U857 ( .A(SRAM_RDATA[1]), .B(MDO[1]), .S(n1980), .Y(
        SRAM_RDATA1309_1) );
    zmux21hb U858 ( .A(SRAM_RDATA[0]), .B(MDO[0]), .S(SRAM_RUN_T), .Y(
        SRAM_RDATA1309_0) );
    zor2b U859 ( .A(WR), .B(WADDR[0]), .Y(WADDR_ATPG1549_0) );
    zor2b U860 ( .A(BIST_RDATA_4), .B(n2019), .Y(BIST_RDATA_T1160_4) );
    zmux21lb U861 ( .A(n2386), .B(n2398), .S(BIST_RDATA_22), .Y(n2139) );
    zmux21lb U862 ( .A(n2404), .B(n2408), .S(BIST_PATTERN[22]), .Y(n2140) );
    zmux21lb U863 ( .A(n2417), .B(n2428), .S(BIST_WDATA_26), .Y(n2079) );
    zmux21lb U864 ( .A(n2438), .B(n1974), .S(BIST_PATTERN[26]), .Y(n2080) );
    zmux21lb U865 ( .A(n2387), .B(n2401), .S(BIST_RDATA_6), .Y(n2106) );
    zmux21lb U866 ( .A(n2285), .B(n2411), .S(BIST_PATTERN[6]), .Y(n2107) );
    zor2b U867 ( .A(BIST_RDATA_12), .B(n2019), .Y(BIST_RDATA_T1160_12) );
    zan2b U868 ( .A(BIST_RDATA_27), .B(n2020), .Y(BIST_RDATA_T1160_27) );
    zmux21lb U869 ( .A(n2414), .B(n2431), .S(BIST_WDATA_2), .Y(n2028) );
    zmux21lb U870 ( .A(n2437), .B(n2443), .S(BIST_PATTERN[2]), .Y(n2029) );
    zmux21lb U871 ( .A(n2421), .B(n2430), .S(BIST_WDATA_13), .Y(n2053) );
    zmux21lb U872 ( .A(n2436), .B(n2442), .S(BIST_PATTERN[13]), .Y(n2054) );
    zmux21lb U873 ( .A(n2285), .B(n2409), .S(BIST_PATTERN[17]), .Y(n2129) );
    zmux21lb U874 ( .A(n2390), .B(n2403), .S(BIST_RDATA_17), .Y(n2130) );
    zmux21lb U875 ( .A(n2390), .B(n2401), .S(BIST_RDATA_30), .Y(n2155) );
    zmux21lb U876 ( .A(n2285), .B(n2411), .S(BIST_PATTERN[30]), .Y(n2156) );
    zmux21lb U877 ( .A(n2288), .B(n2403), .S(BIST_RDATA_10), .Y(n2115) );
    zmux21lb U878 ( .A(n2285), .B(n2412), .S(BIST_PATTERN[10]), .Y(n2116) );
    zmux21lb U879 ( .A(n2421), .B(n2430), .S(BIST_WDATA_28), .Y(n2083) );
    zmux21lb U880 ( .A(n2436), .B(n2442), .S(BIST_PATTERN[28]), .Y(n2084) );
    zmux21lb U881 ( .A(n2391), .B(n2399), .S(BIST_RDATA_8), .Y(n2111) );
    zmux21lb U882 ( .A(n2405), .B(n2409), .S(BIST_PATTERN[8]), .Y(n2112) );
    zmux21lb U883 ( .A(n2420), .B(n2429), .S(BIST_WDATA_14), .Y(n2055) );
    zmux21lb U884 ( .A(n2435), .B(n2441), .S(BIST_PATTERN[14]), .Y(n2056) );
    zmux21lb U885 ( .A(n2415), .B(n2431), .S(BIST_WDATA_5), .Y(n2036) );
    zmux21lb U886 ( .A(n2438), .B(n1974), .S(BIST_PATTERN[5]), .Y(n2037) );
    zor2b U887 ( .A(BIST_RDATA_20), .B(n2019), .Y(BIST_RDATA_T1160_20) );
    zmux21lb U888 ( .A(n2388), .B(n2402), .S(BIST_RDATA_19), .Y(n2133) );
    zmux21lb U889 ( .A(n2406), .B(n1973), .S(BIST_PATTERN[19]), .Y(n2134) );
    zan2b U890 ( .A(BIST_RDATA_15), .B(n2020), .Y(BIST_RDATA_T1160_15) );
    zmux21lb U891 ( .A(n2414), .B(n2429), .S(BIST_WDATA_21), .Y(n2069) );
    zmux21lb U892 ( .A(n2435), .B(n2441), .S(BIST_PATTERN[21]), .Y(n2070) );
    zmux21lb U893 ( .A(n2285), .B(n2412), .S(BIST_PATTERN[1]), .Y(n2094) );
    zmux21lb U894 ( .A(n2288), .B(n2398), .S(BIST_RDATA_1), .Y(n2095) );
    zan2b U895 ( .A(BIST_RDATA_3), .B(n2020), .Y(BIST_RDATA_T1160_3) );
    zan2b U896 ( .A(BIST_RDATA_29), .B(n2020), .Y(BIST_RDATA_T1160_29) );
    zmux21lb U897 ( .A(n2285), .B(n2412), .S(BIST_PATTERN[25]), .Y(n2145) );
    zmux21lb U898 ( .A(n2288), .B(n2403), .S(BIST_RDATA_25), .Y(n2146) );
    zan2b U899 ( .A(BIST_RDATA_21), .B(n2020), .Y(BIST_RDATA_T1160_21) );
    zmux21lb U900 ( .A(n2419), .B(n2428), .S(BIST_WDATA_15), .Y(n2057) );
    zmux21lb U901 ( .A(n2434), .B(n2440), .S(BIST_PATTERN[15]), .Y(n2058) );
    zmux21lb U902 ( .A(n2416), .B(n2432), .S(BIST_WDATA_4), .Y(n2033) );
    zmux21lb U903 ( .A(n2439), .B(n2444), .S(BIST_PATTERN[4]), .Y(n2034) );
    zan2b U904 ( .A(n1950), .B(n2014), .Y(BIST_RUN_C346) );
    zmux21lb U905 ( .A(n2420), .B(n2429), .S(BIST_WDATA_29), .Y(n2085) );
    zmux21lb U906 ( .A(n2435), .B(n2441), .S(BIST_PATTERN[29]), .Y(n2086) );
    zivb U907 ( .A(n2172), .Y(n2379) );
    zivb U908 ( .A(n2169), .Y(n2383) );
    zmux21lb U909 ( .A(n2404), .B(n2408), .S(BIST_PATTERN[9]), .Y(n2113) );
    zmux21lb U910 ( .A(n2386), .B(n2398), .S(BIST_RDATA_9), .Y(n2114) );
    zmux21lb U911 ( .A(n2389), .B(n2402), .S(BIST_RDATA_11), .Y(n2117) );
    zmux21lb U912 ( .A(n2404), .B(n1973), .S(BIST_PATTERN[11]), .Y(n2118) );
    zor2b U913 ( .A(BIST_RDATA_2), .B(n2019), .Y(BIST_RDATA_T1160_2) );
    zor2b U914 ( .A(BIST_RDATA_28), .B(n2019), .Y(BIST_RDATA_T1160_28) );
    zan2b U915 ( .A(n1979), .B(n2013), .Y(SRAM_R_T1481) );
    zivb U916 ( .A(SRAM_WR), .Y(n2013) );
    zmux21lb U917 ( .A(n2288), .B(n2399), .S(BIST_RDATA_24), .Y(n2143) );
    zmux21lb U918 ( .A(n2285), .B(n2412), .S(BIST_PATTERN[24]), .Y(n2144) );
    zmux21lb U919 ( .A(n2416), .B(n2430), .S(BIST_WDATA_20), .Y(n2067) );
    zmux21lb U920 ( .A(n2436), .B(n2442), .S(BIST_PATTERN[20]), .Y(n2068) );
    zmux21lb U921 ( .A(n2288), .B(n2402), .S(BIST_RDATA_0), .Y(n2091) );
    zmux21lb U922 ( .A(n2285), .B(n2408), .S(BIST_PATTERN[0]), .Y(n2092) );
    zmux21lb U923 ( .A(n2389), .B(n2403), .S(BIST_RDATA_18), .Y(n2131) );
    zmux21lb U924 ( .A(n2285), .B(n2412), .S(BIST_PATTERN[18]), .Y(n2132) );
    zor2b U925 ( .A(BIST_RDATA_14), .B(n2019), .Y(BIST_RDATA_T1160_14) );
    zan2b U926 ( .A(BIST_RDATA_13), .B(n2020), .Y(BIST_RDATA_T1160_13) );
    zmux21lb U927 ( .A(n2422), .B(n2431), .S(BIST_WDATA_27), .Y(n2081) );
    zmux21lb U928 ( .A(n2437), .B(n2443), .S(BIST_PATTERN[27]), .Y(n2082) );
    zmux21lb U929 ( .A(n2387), .B(n2400), .S(BIST_RDATA_7), .Y(n2109) );
    zmux21lb U930 ( .A(n2406), .B(n2410), .S(BIST_PATTERN[7]), .Y(n2110) );
    zan2b U931 ( .A(BIST_RDATA_5), .B(n2020), .Y(BIST_RDATA_T1160_5) );
    zmux21lb U932 ( .A(n2288), .B(n2399), .S(BIST_RDATA_23), .Y(n2141) );
    zmux21lb U933 ( .A(n2285), .B(n1973), .S(BIST_PATTERN[23]), .Y(n2142) );
    zmux21lb U934 ( .A(n2390), .B(n2400), .S(BIST_RDATA_16), .Y(n2127) );
    zmux21lb U935 ( .A(n2285), .B(n2410), .S(BIST_PATTERN[16]), .Y(n2128) );
    zor2b U936 ( .A(n2260), .B(n2261), .Y(n2093) );
    zmux21lb U937 ( .A(n2390), .B(n2403), .S(BIST_RDATA_31), .Y(n2157) );
    zmux21lb U938 ( .A(n2285), .B(n2409), .S(BIST_PATTERN[31]), .Y(n2158) );
    zmux21lb U939 ( .A(n2422), .B(n2431), .S(BIST_WDATA_12), .Y(n2051) );
    zmux21lb U940 ( .A(n2437), .B(n2443), .S(BIST_PATTERN[12]), .Y(n2052) );
    zor2b U941 ( .A(n2242), .B(n2245), .Y(n2035) );
    zmux21lb U942 ( .A(n2419), .B(n2428), .S(BIST_WDATA_3), .Y(n2031) );
    zmux21lb U943 ( .A(n2434), .B(n2440), .S(BIST_PATTERN[3]), .Y(n2032) );
    zor2b U944 ( .A(BIST_RDATA_26), .B(n2019), .Y(BIST_RDATA_T1160_26) );
    zmux21lb U945 ( .A(n2288), .B(n2399), .S(BIST_RDATA_21), .Y(n2137) );
    zmux21lb U946 ( .A(n2405), .B(n2409), .S(BIST_PATTERN[21]), .Y(n2138) );
    zan2b U947 ( .A(BIST_RDATA_7), .B(n2020), .Y(BIST_RDATA_T1160_7) );
    zmux21lb U948 ( .A(n2415), .B(n2428), .S(BIST_WDATA_19), .Y(n2065) );
    zmux21lb U949 ( .A(n2438), .B(n1974), .S(BIST_PATTERN[19]), .Y(n2066) );
    zmux21lb U950 ( .A(n2414), .B(n2429), .S(BIST_WDATA_8), .Y(n2043) );
    zmux21lb U951 ( .A(n2435), .B(n2441), .S(BIST_PATTERN[8]), .Y(n2044) );
    zmux21lb U952 ( .A(n2388), .B(n2402), .S(BIST_RDATA_5), .Y(n2104) );
    zmux21lb U953 ( .A(n2406), .B(n1973), .S(BIST_PATTERN[5]), .Y(n2105) );
    zmux21lb U954 ( .A(n2421), .B(n2432), .S(BIST_WDATA_25), .Y(n2077) );
    zmux21lb U955 ( .A(n2439), .B(n2444), .S(BIST_PATTERN[25]), .Y(n2078) );
    zan2b U956 ( .A(BIST_RDATA_11), .B(n2020), .Y(BIST_RDATA_T1160_11) );
    zan2b U957 ( .A(n1736), .B(n2012), .Y(BIST_WR1405) );
    zivb U958 ( .A(n2224), .Y(n2021) );
    zao32b U959 ( .A(n2014), .B(n2015), .C(BIST_WUNDER), .D(BIST_WFULL), .E(
        BISTSM_5), .Y(BIST_RD_T1359) );
    zivb U960 ( .A(n2179), .Y(BIST_WUNDER) );
    zivb U961 ( .A(n2014), .Y(n2377) );
    zivb U962 ( .A(n2015), .Y(BIST_RUNDER) );
    zmux21lb U963 ( .A(n2392), .B(n2400), .S(BIST_RDATA_28), .Y(n2151) );
    zmux21lb U964 ( .A(n2406), .B(n2410), .S(BIST_PATTERN[28]), .Y(n2152) );
    zor2b U965 ( .A(BIST_RDATA_24), .B(n2019), .Y(BIST_RDATA_T1160_24) );
    zmux21lb U966 ( .A(n2420), .B(n2432), .S(BIST_WDATA_1), .Y(n2026) );
    zmux21lb U967 ( .A(n2434), .B(n2444), .S(BIST_PATTERN[1]), .Y(n2027) );
    zmux21lb U968 ( .A(n2422), .B(n2432), .S(BIST_WDATA_10), .Y(n2047) );
    zmux21lb U969 ( .A(n2439), .B(n2444), .S(BIST_PATTERN[10]), .Y(n2048) );
    zor2b U970 ( .A(BIST_RDATA_18), .B(n2019), .Y(BIST_RDATA_T1160_18) );
    zan2b U971 ( .A(SRAM_WR), .B(n1978), .Y(SRAM_W_T1443) );
    zmux21lb U972 ( .A(n2391), .B(n2399), .S(BIST_RDATA_14), .Y(n2123) );
    zmux21lb U973 ( .A(n2405), .B(n2409), .S(BIST_PATTERN[14]), .Y(n2124) );
    zor2b U974 ( .A(n2260), .B(n2262), .Y(n2108) );
    zmux21lb U975 ( .A(n2392), .B(n2400), .S(BIST_RDATA_13), .Y(n2121) );
    zmux21lb U976 ( .A(n2406), .B(n2410), .S(BIST_PATTERN[13]), .Y(n2122) );
    zmux21lb U977 ( .A(n2418), .B(n2431), .S(BIST_WDATA_30), .Y(n2087) );
    zmux21lb U978 ( .A(n2439), .B(n2443), .S(BIST_PATTERN[30]), .Y(n2088) );
    zmux21lb U979 ( .A(n2417), .B(n2429), .S(BIST_WDATA_17), .Y(n2061) );
    zmux21lb U980 ( .A(n2438), .B(n2441), .S(BIST_PATTERN[17]), .Y(n2062) );
    zmux21lb U981 ( .A(n2413), .B(n2431), .S(BIST_WDATA_6), .Y(n2038) );
    zmux21lb U982 ( .A(n2437), .B(n2443), .S(BIST_PATTERN[6]), .Y(n2039) );
    zan2b U983 ( .A(BIST_RDATA_9), .B(n2020), .Y(BIST_RDATA_T1160_9) );
    zan2b U984 ( .A(BIST_RDATA_23), .B(n2020), .Y(BIST_RDATA_T1160_23) );
    zan2b U985 ( .A(BIST_RDATA_31), .B(n2020), .Y(BIST_RDATA_T1160_31) );
    zor2b U986 ( .A(BIST_RDATA_16), .B(n2019), .Y(BIST_RDATA_T1160_16) );
    zmux21lb U987 ( .A(n2413), .B(n2428), .S(BIST_WDATA_22), .Y(n2071) );
    zmux21lb U988 ( .A(n2434), .B(n2440), .S(BIST_PATTERN[22]), .Y(n2072) );
    zor2b U989 ( .A(n2242), .B(n2244), .Y(n2040) );
    zmux21lb U990 ( .A(n2386), .B(n2401), .S(BIST_RDATA_2), .Y(n2096) );
    zmux21lb U991 ( .A(n2404), .B(n2411), .S(BIST_PATTERN[2]), .Y(n2097) );
    zmux21lb U992 ( .A(n2391), .B(n2402), .S(BIST_RDATA_26), .Y(n2147) );
    zmux21lb U993 ( .A(n2405), .B(n1973), .S(BIST_PATTERN[26]), .Y(n2148) );
    zor2b U994 ( .A(n2260), .B(n2264), .Y(n2098) );
    zor2b U995 ( .A(BIST_RDATA_0), .B(n2019), .Y(BIST_RDATA_T1160_0) );
    zor2b U996 ( .A(BIST_RDATA_8), .B(n2019), .Y(BIST_RDATA_T1160_8) );
    zor2b U997 ( .A(BIST_RDATA_22), .B(n2019), .Y(BIST_RDATA_T1160_22) );
    zmux21lb U998 ( .A(n2417), .B(n2429), .S(BIST_WDATA_31), .Y(n2089) );
    zmux21lb U999 ( .A(n2435), .B(n2441), .S(BIST_PATTERN[31]), .Y(n2090) );
    zmux21lb U1000 ( .A(n2418), .B(n2430), .S(BIST_WDATA_16), .Y(n2059) );
    zmux21lb U1001 ( .A(n2437), .B(n2442), .S(BIST_PATTERN[16]), .Y(n2060) );
    zmux21lb U1002 ( .A(n2422), .B(n2430), .S(BIST_WDATA_7), .Y(n2041) );
    zmux21lb U1003 ( .A(n2436), .B(n2442), .S(BIST_PATTERN[7]), .Y(n2042) );
    zmux21lb U1004 ( .A(n2392), .B(n2401), .S(BIST_RDATA_12), .Y(n2119) );
    zmux21lb U1005 ( .A(n2285), .B(n2411), .S(BIST_PATTERN[12]), .Y(n2120) );
    zmux21lb U1006 ( .A(n2392), .B(n2401), .S(BIST_RDATA_27), .Y(n2149) );
    zmux21lb U1007 ( .A(n2285), .B(n2411), .S(BIST_PATTERN[27]), .Y(n2150) );
    zan2b U1008 ( .A(BIST_RDATA_1), .B(n2020), .Y(BIST_RDATA_T1160_1) );
    zmux21lb U1009 ( .A(n2388), .B(n2398), .S(BIST_RDATA_3), .Y(n2099) );
    zmux21lb U1010 ( .A(n2404), .B(n2408), .S(BIST_PATTERN[3]), .Y(n2100) );
    zivb U1011 ( .A(n2167), .Y(n2385) );
    zan2b U1012 ( .A(SLREAD), .B(SLAVEMODE), .Y(RPOP187) );
    zmux21lb U1013 ( .A(n2416), .B(n2430), .S(BIST_WDATA_23), .Y(n2073) );
    zmux21lb U1014 ( .A(n2436), .B(n1974), .S(BIST_PATTERN[23]), .Y(n2074) );
    zor2b U1015 ( .A(BIST_RDATA_30), .B(n2019), .Y(BIST_RDATA_T1160_30) );
    zan2b U1016 ( .A(BIST_RDATA_17), .B(n2020), .Y(BIST_RDATA_T1160_17) );
    zao32b U1017 ( .A(n2016), .B(n2009), .C(BIST_WFULL), .D(n2017), .E(
        BIST_RD_T), .Y(BIST_RD1353) );
    zivb U1018 ( .A(n2236), .Y(BIST_WFULL) );
    znd8b U1019 ( .A(n2215), .B(n2216), .C(n2217), .D(n2218), .E(n2183), .F(
        n2184), .G(BIST_WADDR_0), .H(n2255), .Y(n2236) );
    zivb U1020 ( .A(n2009), .Y(BIST_RFULL) );
    zor2b U1021 ( .A(BIST_RDATA_10), .B(n2019), .Y(BIST_RDATA_T1160_10) );
    zmux21lb U1022 ( .A(n2419), .B(n2432), .S(BIST_WDATA_24), .Y(n2075) );
    zmux21lb U1023 ( .A(n2435), .B(n2444), .S(BIST_PATTERN[24]), .Y(n2076) );
    zmux21lb U1024 ( .A(n2389), .B(n2403), .S(BIST_RDATA_4), .Y(n2101) );
    zmux21lb U1025 ( .A(n2285), .B(n2412), .S(BIST_PATTERN[4]), .Y(n2102) );
    zmux21lb U1026 ( .A(n2416), .B(n2432), .S(BIST_WDATA_18), .Y(n2063) );
    zmux21lb U1027 ( .A(n2439), .B(n2444), .S(BIST_PATTERN[18]), .Y(n2064) );
    zor2b U1028 ( .A(n2242), .B(n2246), .Y(n2030) );
    zmux21lb U1029 ( .A(n2413), .B(n2428), .S(BIST_WDATA_9), .Y(n2045) );
    zmux21lb U1030 ( .A(n2434), .B(n2440), .S(BIST_PATTERN[9]), .Y(n2046) );
    zivb U1031 ( .A(n2176), .Y(n2378) );
    zmux21lb U1032 ( .A(n2387), .B(n2400), .S(BIST_RDATA_20), .Y(n2135) );
    zmux21lb U1033 ( .A(n2406), .B(n2410), .S(BIST_PATTERN[20]), .Y(n2136) );
    zor2b U1034 ( .A(n2260), .B(n2263), .Y(n2103) );
    zivb U1035 ( .A(n2374), .Y(n2260) );
    zor2b U1036 ( .A(BIST_RDATA_6), .B(n2019), .Y(BIST_RDATA_T1160_6) );
    zan2b U1037 ( .A(BIST_RDATA_19), .B(n2020), .Y(BIST_RDATA_T1160_19) );
    zmux21lb U1038 ( .A(n2388), .B(n2398), .S(BIST_RDATA_15), .Y(n2125) );
    zmux21lb U1039 ( .A(n2404), .B(n2408), .S(BIST_PATTERN[15]), .Y(n2126) );
    zmux21lb U1040 ( .A(n2418), .B(n2430), .S(BIST_WDATA_11), .Y(n2049) );
    zmux21lb U1041 ( .A(n2438), .B(n1974), .S(BIST_PATTERN[11]), .Y(n2050) );
    zivb U1042 ( .A(n2277), .Y(n2369) );
    zivb U1043 ( .A(n2174), .Y(n2380) );
    zmux21lb U1044 ( .A(n2415), .B(n2428), .S(BIST_WDATA_0), .Y(n2023) );
    zmux21lb U1045 ( .A(n2434), .B(n2440), .S(BIST_PATTERN[0]), .Y(n2024) );
    zor2b U1046 ( .A(n2242), .B(n2243), .Y(n2025) );
    zivb U1047 ( .A(n2370), .Y(n2242) );
    zmux21lb U1048 ( .A(n2391), .B(n2399), .S(BIST_RDATA_29), .Y(n2153) );
    zmux21lb U1049 ( .A(n2405), .B(n2409), .S(BIST_PATTERN[29]), .Y(n2154) );
    zivb U1050 ( .A(n2290), .Y(n2373) );
    zivb U1051 ( .A(n2291), .Y(n2381) );
    zivb U1052 ( .A(n2165), .Y(n2384) );
    zan2b U1053 ( .A(BIST_RDATA_25), .B(n2020), .Y(BIST_RDATA_T1160_25) );
    zivb U1054 ( .A(n2196), .Y(BISTSMNXT_5) );
    zivb U1055 ( .A(n2020), .Y(n2019) );
    zmux31hb U1056 ( .A(n1975), .B(n1976), .D0(WMA[0]), .D1(SRAM_ADDR[0]), 
        .D2(BIST_WADDR_0), .Y(WADDR[0]) );
    zmux31hb U1057 ( .A(n1978), .B(n1976), .D0(WMA[1]), .D1(SRAM_ADDR[1]), 
        .D2(BIST_WADDR_1), .Y(WADDR[1]) );
    zmux31hb U1058 ( .A(n1979), .B(n1972), .D0(WMA[2]), .D1(SRAM_ADDR[2]), 
        .D2(BIST_WADDR_2), .Y(WADDR[2]) );
    zmux31hb U1059 ( .A(n1979), .B(n1972), .D0(WMA[3]), .D1(SRAM_ADDR[3]), 
        .D2(BIST_WADDR_3), .Y(WADDR[3]) );
    zmux31hb U1060 ( .A(n1978), .B(n1976), .D0(WMA[4]), .D1(SRAM_ADDR[4]), 
        .D2(BIST_WADDR_4), .Y(WADDR[4]) );
    zmux31hb U1061 ( .A(n1979), .B(n1976), .D0(WMA[5]), .D1(SRAM_ADDR[5]), 
        .D2(BIST_WADDR_5), .Y(WADDR[5]) );
    zmux31hb U1062 ( .A(n1978), .B(n1976), .D0(WMA[6]), .D1(SRAM_ADDR[6]), 
        .D2(BIST_WADDR_6), .Y(WADDR[6]) );
    zmux31hb U1063 ( .A(n1975), .B(n1976), .D0(WMA[7]), .D1(SRAM_ADDR[7]), 
        .D2(BIST_WADDR_7), .Y(WADDR[7]) );
    zmux31hb U1064 ( .A(n1979), .B(n1976), .D0(WMA[8]), .D1(SRAM_ADDR[8]), 
        .D2(BIST_WADDR_8), .Y(WADDR[8]) );
    zmux31hb U1065 ( .A(n1978), .B(n1740), .D0(FIFO_MDI[0]), .D1(BIST_PATTERN
        [0]), .D2(BIST_WDATA_0), .Y(MDI[0]) );
    zmux31hb U1066 ( .A(n1975), .B(n1740), .D0(FIFO_MDI[1]), .D1(BIST_PATTERN
        [1]), .D2(BIST_WDATA_1), .Y(MDI[1]) );
    zmux31hb U1067 ( .A(n1979), .B(n1976), .D0(FIFO_MDI[2]), .D1(BIST_PATTERN
        [2]), .D2(BIST_WDATA_2), .Y(MDI[2]) );
    zmux31hb U1068 ( .A(n1979), .B(n1740), .D0(FIFO_MDI[3]), .D1(BIST_PATTERN
        [3]), .D2(BIST_WDATA_3), .Y(MDI[3]) );
    zmux31hb U1069 ( .A(n1975), .B(n1740), .D0(FIFO_MDI[4]), .D1(BIST_PATTERN
        [4]), .D2(BIST_WDATA_4), .Y(MDI[4]) );
    zmux31hb U1070 ( .A(n1975), .B(n1976), .D0(FIFO_MDI[5]), .D1(BIST_PATTERN
        [5]), .D2(BIST_WDATA_5), .Y(MDI[5]) );
    zmux31hb U1071 ( .A(n1979), .B(n1740), .D0(FIFO_MDI[6]), .D1(BIST_PATTERN
        [6]), .D2(BIST_WDATA_6), .Y(MDI[6]) );
    zmux31hb U1072 ( .A(n1978), .B(n1740), .D0(FIFO_MDI[7]), .D1(BIST_PATTERN
        [7]), .D2(BIST_WDATA_7), .Y(MDI[7]) );
    zmux31hb U1073 ( .A(n1979), .B(n1740), .D0(FIFO_MDI[8]), .D1(BIST_PATTERN
        [8]), .D2(BIST_WDATA_8), .Y(MDI[8]) );
    zmux31hb U1074 ( .A(n1978), .B(n1740), .D0(FIFO_MDI[9]), .D1(BIST_PATTERN
        [9]), .D2(BIST_WDATA_9), .Y(MDI[9]) );
    zmux31hb U1075 ( .A(n1979), .B(n1740), .D0(FIFO_MDI[10]), .D1(BIST_PATTERN
        [10]), .D2(BIST_WDATA_10), .Y(MDI[10]) );
    zmux31hb U1076 ( .A(n1979), .B(n1976), .D0(FIFO_MDI[11]), .D1(BIST_PATTERN
        [11]), .D2(BIST_WDATA_11), .Y(MDI[11]) );
    zmux31hb U1077 ( .A(n1975), .B(n1976), .D0(FIFO_MDI[12]), .D1(BIST_PATTERN
        [12]), .D2(BIST_WDATA_12), .Y(MDI[12]) );
    zmux31hb U1078 ( .A(n1978), .B(n1972), .D0(FIFO_MDI[13]), .D1(BIST_PATTERN
        [13]), .D2(BIST_WDATA_13), .Y(MDI[13]) );
    zmux31hb U1079 ( .A(n1978), .B(n1740), .D0(FIFO_MDI[14]), .D1(BIST_PATTERN
        [14]), .D2(BIST_WDATA_14), .Y(MDI[14]) );
    zmux31hb U1080 ( .A(n1975), .B(n1740), .D0(FIFO_MDI[15]), .D1(BIST_PATTERN
        [15]), .D2(BIST_WDATA_15), .Y(MDI[15]) );
    zmux31hb U1081 ( .A(n1978), .B(n1740), .D0(FIFO_MDI[16]), .D1(BIST_PATTERN
        [16]), .D2(BIST_WDATA_16), .Y(MDI[16]) );
    zmux31hb U1082 ( .A(n1975), .B(n1976), .D0(FIFO_MDI[17]), .D1(BIST_PATTERN
        [17]), .D2(BIST_WDATA_17), .Y(MDI[17]) );
    zmux31hb U1083 ( .A(n1975), .B(n1976), .D0(FIFO_MDI[18]), .D1(BIST_PATTERN
        [18]), .D2(BIST_WDATA_18), .Y(MDI[18]) );
    zmux31hb U1084 ( .A(n1979), .B(n1740), .D0(FIFO_MDI[19]), .D1(BIST_PATTERN
        [19]), .D2(BIST_WDATA_19), .Y(MDI[19]) );
    zmux31hb U1085 ( .A(n1979), .B(n1740), .D0(FIFO_MDI[20]), .D1(BIST_PATTERN
        [20]), .D2(BIST_WDATA_20), .Y(MDI[20]) );
    zmux31hb U1086 ( .A(n1978), .B(n1976), .D0(FIFO_MDI[21]), .D1(BIST_PATTERN
        [21]), .D2(BIST_WDATA_21), .Y(MDI[21]) );
    zmux31hb U1087 ( .A(n1975), .B(n1740), .D0(FIFO_MDI[22]), .D1(BIST_PATTERN
        [22]), .D2(BIST_WDATA_22), .Y(MDI[22]) );
    zmux31hb U1088 ( .A(n1975), .B(n1976), .D0(FIFO_MDI[23]), .D1(BIST_PATTERN
        [23]), .D2(BIST_WDATA_23), .Y(MDI[23]) );
    zmux31hb U1089 ( .A(n1975), .B(n1976), .D0(FIFO_MDI[24]), .D1(BIST_PATTERN
        [24]), .D2(BIST_WDATA_24), .Y(MDI[24]) );
    zmux31hb U1090 ( .A(n1978), .B(n1976), .D0(FIFO_MDI[25]), .D1(BIST_PATTERN
        [25]), .D2(BIST_WDATA_25), .Y(MDI[25]) );
    zmux31hb U1091 ( .A(n1978), .B(n1976), .D0(FIFO_MDI[26]), .D1(BIST_PATTERN
        [26]), .D2(BIST_WDATA_26), .Y(MDI[26]) );
    zmux31hb U1092 ( .A(n1975), .B(n1740), .D0(FIFO_MDI[27]), .D1(BIST_PATTERN
        [27]), .D2(BIST_WDATA_27), .Y(MDI[27]) );
    zmux31hb U1093 ( .A(n1975), .B(n1976), .D0(FIFO_MDI[28]), .D1(BIST_PATTERN
        [28]), .D2(BIST_WDATA_28), .Y(MDI[28]) );
    zmux31hb U1094 ( .A(n1979), .B(n1740), .D0(FIFO_MDI[29]), .D1(BIST_PATTERN
        [29]), .D2(BIST_WDATA_29), .Y(MDI[29]) );
    zmux31hb U1095 ( .A(n1978), .B(n1740), .D0(FIFO_MDI[30]), .D1(BIST_PATTERN
        [30]), .D2(BIST_WDATA_30), .Y(MDI[30]) );
    zmux31hb U1096 ( .A(n1979), .B(n1740), .D0(FIFO_MDI[31]), .D1(BIST_PATTERN
        [31]), .D2(BIST_WDATA_31), .Y(MDI[31]) );
    zivc U1097 ( .A(n1971), .Y(n1740) );
    zmux21hb U1098 ( .A(n2265), .B(RPOP), .S(SLAVEMODE), .Y(RD) );
    zmux31lb U1099 ( .A(SLAVEMODE), .B(n1979), .D0(n2007), .D1(n2006), .D2(
        n2005), .Y(RADDR[0]) );
    zmux21lb U1100 ( .A(RMA[0]), .B(BIST_RADDR_0), .S(n1736), .Y(n2007) );
    zmux21lb U1101 ( .A(SLADDR[0]), .B(BIST_RADDR_0), .S(n1972), .Y(n2006) );
    zmux21lb U1102 ( .A(SRAM_ADDR[0]), .B(BIST_RADDR_0), .S(n1972), .Y(n2005)
         );
    zmux31lb U1103 ( .A(SLAVEMODE), .B(n1979), .D0(n2004), .D1(n2003), .D2(
        n2002), .Y(RADDR[1]) );
    zmux21lb U1104 ( .A(RMA[1]), .B(BIST_RADDR_1), .S(n1972), .Y(n2004) );
    zmux21lb U1105 ( .A(SLADDR[1]), .B(BIST_RADDR_1), .S(n1972), .Y(n2003) );
    zmux21lb U1106 ( .A(SRAM_ADDR[1]), .B(BIST_RADDR_1), .S(n1972), .Y(n2002)
         );
    zmux31lb U1107 ( .A(SLAVEMODE), .B(n1975), .D0(n2001), .D1(n2000), .D2(
        n1999), .Y(RADDR[2]) );
    zmux21lb U1108 ( .A(RMA[2]), .B(BIST_RADDR_2), .S(n1736), .Y(n2001) );
    zmux21lb U1109 ( .A(SLADDR[2]), .B(BIST_RADDR_2), .S(n1736), .Y(n2000) );
    zmux21lb U1110 ( .A(SRAM_ADDR[2]), .B(BIST_RADDR_2), .S(n1972), .Y(n1999)
         );
    zmux31lb U1111 ( .A(SLAVEMODE), .B(n1978), .D0(n1998), .D1(n1997), .D2(
        n1996), .Y(RADDR[3]) );
    zmux21lb U1112 ( .A(RMA[3]), .B(BIST_RADDR_3), .S(n1736), .Y(n1998) );
    zmux21lb U1113 ( .A(SLADDR[3]), .B(BIST_RADDR_3), .S(n1972), .Y(n1997) );
    zmux21lb U1114 ( .A(SRAM_ADDR[3]), .B(BIST_RADDR_3), .S(n1736), .Y(n1996)
         );
    zmux31lb U1115 ( .A(SLAVEMODE), .B(n1978), .D0(n1995), .D1(n1994), .D2(
        n1993), .Y(RADDR[4]) );
    zmux21lb U1116 ( .A(RMA[4]), .B(BIST_RADDR_4), .S(n1972), .Y(n1995) );
    zmux21lb U1117 ( .A(SLADDR[4]), .B(BIST_RADDR_4), .S(n1736), .Y(n1994) );
    zmux21lb U1118 ( .A(SRAM_ADDR[4]), .B(BIST_RADDR_4), .S(n1972), .Y(n1993)
         );
    zmux31lb U1119 ( .A(SLAVEMODE), .B(n1978), .D0(n1992), .D1(n1991), .D2(
        n1990), .Y(RADDR[5]) );
    zmux21lb U1120 ( .A(RMA[5]), .B(BIST_RADDR_5), .S(n1736), .Y(n1992) );
    zmux21lb U1121 ( .A(SLADDR[5]), .B(BIST_RADDR_5), .S(n1972), .Y(n1991) );
    zmux21lb U1122 ( .A(SRAM_ADDR[5]), .B(BIST_RADDR_5), .S(n1972), .Y(n1990)
         );
    zmux31lb U1123 ( .A(SLAVEMODE), .B(n1979), .D0(n1989), .D1(n1988), .D2(
        n1987), .Y(RADDR[6]) );
    zmux21lb U1124 ( .A(RMA[6]), .B(BIST_RADDR_6), .S(n1972), .Y(n1989) );
    zmux21lb U1125 ( .A(SLADDR[6]), .B(BIST_RADDR_6), .S(n1736), .Y(n1988) );
    zmux21lb U1126 ( .A(SRAM_ADDR[6]), .B(BIST_RADDR_6), .S(n1736), .Y(n1987)
         );
    zmux31lb U1127 ( .A(SLAVEMODE), .B(n1975), .D0(n1986), .D1(n1985), .D2(
        n1984), .Y(RADDR[7]) );
    zmux21lb U1128 ( .A(RMA[7]), .B(BIST_RADDR_7), .S(n1972), .Y(n1986) );
    zmux21lb U1129 ( .A(SLADDR[7]), .B(BIST_RADDR_7), .S(n1736), .Y(n1985) );
    zmux21lb U1130 ( .A(SRAM_ADDR[7]), .B(BIST_RADDR_7), .S(n1972), .Y(n1984)
         );
    zmux21lb U1131 ( .A(n1982), .B(n1981), .S(n1978), .Y(RADDR[8]) );
    zmux21lb U1132 ( .A(n1983), .B(BIST_RADDR_8), .S(n1972), .Y(n1982) );
    zmux21lb U1133 ( .A(SRAM_ADDR[8]), .B(BIST_RADDR_8), .S(n1736), .Y(n1981)
         );
    zdffqrb BISTSM_reg_8 ( .CK(PCICLK), .D(n1950), .R(TRST_), .Q(BISTSM_8) );
    zivb U1134 ( .A(BISTSM_8), .Y(n2206) );
    zdffqrb BISTSM_reg_7 ( .CK(PCICLK), .D(BISTSMNXT_7), .R(TRST_), .Q(
        BISTSM_7) );
    zdffqrb BISTSM_reg_6 ( .CK(PCICLK), .D(BISTSMNXT_6), .R(TRST_), .Q(
        BISTSM_6) );
    zivb U1135 ( .A(BISTSM_6), .Y(n2227) );
    zdffqrb BISTSM_reg_5 ( .CK(PCICLK), .D(BISTSMNXT_5), .R(TRST_), .Q(
        BISTSM_5) );
    zivb U1136 ( .A(BISTSM_5), .Y(n2228) );
    zdffqrb BISTSM_reg_4 ( .CK(PCICLK), .D(BISTSMNXT_4), .R(TRST_), .Q(
        BISTSM_4) );
    zivb U1137 ( .A(BISTSM_4), .Y(n2222) );
    zdffqrb BISTSM_reg_3 ( .CK(PCICLK), .D(BISTSMNXT_3), .R(TRST_), .Q(
        BISTSM_3) );
    zivb U1138 ( .A(BISTSM_3), .Y(n2226) );
    zdffqrb BISTSM_reg_2 ( .CK(PCICLK), .D(BISTSMNXT_2), .R(TRST_), .Q(
        BISTSM_2) );
    zivb U1139 ( .A(BISTSM_2), .Y(n2232) );
    zdffrb BISTSM_reg_1 ( .CK(PCICLK), .D(n1952), .R(TRST_), .Q(BISTSM_1), 
        .QN(n2187) );
    zdffqrb BISTSM_reg_0 ( .CK(PCICLK), .D(n1951), .R(TRST_), .Q(BISTSM_0) );
    zivb U1140 ( .A(BISTSM_0), .Y(n2234) );
    zdffqrb BIST_WADDR_reg_8 ( .CK(PCICLK), .D(BIST_WADDR677_8), .R(TRST_), 
        .Q(BIST_WADDR_8) );
    zivb U1141 ( .A(BIST_WADDR_8), .Y(n2181) );
    zdffqrb BIST_WADDR_reg_7 ( .CK(PCICLK), .D(BIST_WADDR677_7), .R(TRST_), 
        .Q(BIST_WADDR_7) );
    zivb U1142 ( .A(BIST_WADDR_7), .Y(n2182) );
    zdffqrb BIST_WADDR_reg_6 ( .CK(PCICLK), .D(BIST_WADDR677_6), .R(TRST_), 
        .Q(BIST_WADDR_6) );
    zivb U1143 ( .A(BIST_WADDR_6), .Y(n2218) );
    zdffqrb BIST_WADDR_reg_5 ( .CK(PCICLK), .D(BIST_WADDR677_5), .R(TRST_), 
        .Q(BIST_WADDR_5) );
    zivb U1144 ( .A(BIST_WADDR_5), .Y(n2217) );
    zdffqrb BIST_WADDR_reg_4 ( .CK(PCICLK), .D(BIST_WADDR677_4), .R(TRST_), 
        .Q(BIST_WADDR_4) );
    zivb U1145 ( .A(BIST_WADDR_4), .Y(n2216) );
    zdffqrb BIST_WADDR_reg_3 ( .CK(PCICLK), .D(BIST_WADDR677_3), .R(TRST_), 
        .Q(BIST_WADDR_3) );
    zivb U1146 ( .A(BIST_WADDR_3), .Y(n2215) );
    zdffqrb BIST_WADDR_reg_2 ( .CK(PCICLK), .D(BIST_WADDR677_2), .R(TRST_), 
        .Q(BIST_WADDR_2) );
    zivb U1147 ( .A(BIST_WADDR_2), .Y(n2184) );
    zdffqrb BIST_WADDR_reg_1 ( .CK(PCICLK), .D(BIST_WADDR677_1), .R(TRST_), 
        .Q(BIST_WADDR_1) );
    zivb U1148 ( .A(BIST_WADDR_1), .Y(n2183) );
    zdffqrb BIST_WADDR_reg_0 ( .CK(PCICLK), .D(BIST_WADDR677_0), .R(TRST_), 
        .Q(BIST_WADDR_0) );
    zivb U1149 ( .A(BIST_WADDR_0), .Y(n2180) );
    zdffqrb BIST_RADDR_reg_8 ( .CK(PCICLK), .D(BIST_RADDR1065_8), .R(TRST_), 
        .Q(BIST_RADDR_8) );
    zivb U1150 ( .A(BIST_RADDR_8), .Y(n2200) );
    zdffqrb BIST_RADDR_reg_7 ( .CK(PCICLK), .D(BIST_RADDR1065_7), .R(TRST_), 
        .Q(BIST_RADDR_7) );
    zivb U1151 ( .A(BIST_RADDR_7), .Y(n2203) );
    zdffqrb BIST_RADDR_reg_6 ( .CK(PCICLK), .D(BIST_RADDR1065_6), .R(TRST_), 
        .Q(BIST_RADDR_6) );
    zivb U1152 ( .A(BIST_RADDR_6), .Y(n2254) );
    zdffqrb BIST_RADDR_reg_5 ( .CK(PCICLK), .D(BIST_RADDR1065_5), .R(TRST_), 
        .Q(BIST_RADDR_5) );
    zivb U1153 ( .A(BIST_RADDR_5), .Y(n2253) );
    zdffqrb BIST_RADDR_reg_4 ( .CK(PCICLK), .D(BIST_RADDR1065_4), .R(TRST_), 
        .Q(BIST_RADDR_4) );
    zivb U1154 ( .A(BIST_RADDR_4), .Y(n2252) );
    zdffqrb BIST_RADDR_reg_3 ( .CK(PCICLK), .D(BIST_RADDR1065_3), .R(TRST_), 
        .Q(BIST_RADDR_3) );
    zivb U1155 ( .A(BIST_RADDR_3), .Y(n2251) );
    zdffqrb BIST_RADDR_reg_2 ( .CK(PCICLK), .D(BIST_RADDR1065_2), .R(TRST_), 
        .Q(BIST_RADDR_2) );
    zivb U1156 ( .A(BIST_RADDR_2), .Y(n2250) );
    zdffqrb BIST_RADDR_reg_1 ( .CK(PCICLK), .D(BIST_RADDR1065_1), .R(TRST_), 
        .Q(BIST_RADDR_1) );
    zivb U1157 ( .A(BIST_RADDR_1), .Y(n2249) );
    zdffqrb BIST_RADDR_reg_0 ( .CK(PCICLK), .D(BIST_RADDR1065_0), .R(TRST_), 
        .Q(BIST_RADDR_0) );
    zivb U1158 ( .A(BIST_RADDR_0), .Y(n2220) );
    zdffqrb SRAM_RDATA_reg_31 ( .CK(PCICLK), .D(SRAM_RDATA1309_31), .R(TRST_), 
        .Q(SRAM_RDATA[31]) );
    zdffqrb SRAM_RDATA_reg_30 ( .CK(PCICLK), .D(SRAM_RDATA1309_30), .R(TRST_), 
        .Q(SRAM_RDATA[30]) );
    zdffqrb SRAM_RDATA_reg_29 ( .CK(PCICLK), .D(SRAM_RDATA1309_29), .R(TRST_), 
        .Q(SRAM_RDATA[29]) );
    zdffqrb SRAM_RDATA_reg_28 ( .CK(PCICLK), .D(SRAM_RDATA1309_28), .R(TRST_), 
        .Q(SRAM_RDATA[28]) );
    zdffqrb SRAM_RDATA_reg_27 ( .CK(PCICLK), .D(SRAM_RDATA1309_27), .R(TRST_), 
        .Q(SRAM_RDATA[27]) );
    zdffqrb SRAM_RDATA_reg_26 ( .CK(PCICLK), .D(SRAM_RDATA1309_26), .R(TRST_), 
        .Q(SRAM_RDATA[26]) );
    zdffqrb SRAM_RDATA_reg_25 ( .CK(PCICLK), .D(SRAM_RDATA1309_25), .R(TRST_), 
        .Q(SRAM_RDATA[25]) );
    zdffqrb SRAM_RDATA_reg_24 ( .CK(PCICLK), .D(SRAM_RDATA1309_24), .R(TRST_), 
        .Q(SRAM_RDATA[24]) );
    zdffqrb SRAM_RDATA_reg_23 ( .CK(PCICLK), .D(SRAM_RDATA1309_23), .R(TRST_), 
        .Q(SRAM_RDATA[23]) );
    zdffqrb SRAM_RDATA_reg_22 ( .CK(PCICLK), .D(SRAM_RDATA1309_22), .R(TRST_), 
        .Q(SRAM_RDATA[22]) );
    zdffqrb SRAM_RDATA_reg_21 ( .CK(PCICLK), .D(SRAM_RDATA1309_21), .R(TRST_), 
        .Q(SRAM_RDATA[21]) );
    zdffqrb SRAM_RDATA_reg_20 ( .CK(PCICLK), .D(SRAM_RDATA1309_20), .R(TRST_), 
        .Q(SRAM_RDATA[20]) );
    zdffqrb SRAM_RDATA_reg_19 ( .CK(PCICLK), .D(SRAM_RDATA1309_19), .R(TRST_), 
        .Q(SRAM_RDATA[19]) );
    zdffqrb SRAM_RDATA_reg_18 ( .CK(PCICLK), .D(SRAM_RDATA1309_18), .R(TRST_), 
        .Q(SRAM_RDATA[18]) );
    zdffqrb SRAM_RDATA_reg_17 ( .CK(PCICLK), .D(SRAM_RDATA1309_17), .R(TRST_), 
        .Q(SRAM_RDATA[17]) );
    zdffqrb SRAM_RDATA_reg_16 ( .CK(PCICLK), .D(SRAM_RDATA1309_16), .R(TRST_), 
        .Q(SRAM_RDATA[16]) );
    zdffqrb SRAM_RDATA_reg_15 ( .CK(PCICLK), .D(SRAM_RDATA1309_15), .R(TRST_), 
        .Q(SRAM_RDATA[15]) );
    zdffqrb SRAM_RDATA_reg_14 ( .CK(PCICLK), .D(SRAM_RDATA1309_14), .R(TRST_), 
        .Q(SRAM_RDATA[14]) );
    zdffqrb SRAM_RDATA_reg_13 ( .CK(PCICLK), .D(SRAM_RDATA1309_13), .R(TRST_), 
        .Q(SRAM_RDATA[13]) );
    zdffqrb SRAM_RDATA_reg_12 ( .CK(PCICLK), .D(SRAM_RDATA1309_12), .R(TRST_), 
        .Q(SRAM_RDATA[12]) );
    zdffqrb SRAM_RDATA_reg_11 ( .CK(PCICLK), .D(SRAM_RDATA1309_11), .R(TRST_), 
        .Q(SRAM_RDATA[11]) );
    zdffqrb SRAM_RDATA_reg_10 ( .CK(PCICLK), .D(SRAM_RDATA1309_10), .R(TRST_), 
        .Q(SRAM_RDATA[10]) );
    zdffqrb SRAM_RDATA_reg_9 ( .CK(PCICLK), .D(SRAM_RDATA1309_9), .R(TRST_), 
        .Q(SRAM_RDATA[9]) );
    zdffqrb SRAM_RDATA_reg_8 ( .CK(PCICLK), .D(SRAM_RDATA1309_8), .R(TRST_), 
        .Q(SRAM_RDATA[8]) );
    zdffqrb SRAM_RDATA_reg_7 ( .CK(PCICLK), .D(SRAM_RDATA1309_7), .R(TRST_), 
        .Q(SRAM_RDATA[7]) );
    zdffqrb SRAM_RDATA_reg_6 ( .CK(PCICLK), .D(SRAM_RDATA1309_6), .R(TRST_), 
        .Q(SRAM_RDATA[6]) );
    zdffqrb SRAM_RDATA_reg_5 ( .CK(PCICLK), .D(SRAM_RDATA1309_5), .R(TRST_), 
        .Q(SRAM_RDATA[5]) );
    zdffqrb SRAM_RDATA_reg_4 ( .CK(PCICLK), .D(SRAM_RDATA1309_4), .R(TRST_), 
        .Q(SRAM_RDATA[4]) );
    zdffqrb SRAM_RDATA_reg_3 ( .CK(PCICLK), .D(SRAM_RDATA1309_3), .R(TRST_), 
        .Q(SRAM_RDATA[3]) );
    zdffqrb SRAM_RDATA_reg_2 ( .CK(PCICLK), .D(SRAM_RDATA1309_2), .R(TRST_), 
        .Q(SRAM_RDATA[2]) );
    zdffqrb SRAM_RDATA_reg_1 ( .CK(PCICLK), .D(SRAM_RDATA1309_1), .R(TRST_), 
        .Q(SRAM_RDATA[1]) );
    zdffqrb SRAM_RDATA_reg_0 ( .CK(PCICLK), .D(SRAM_RDATA1309_0), .R(TRST_), 
        .Q(SRAM_RDATA[0]) );
    zdffqsb BIST_RDATA_T_reg_4 ( .CK(PCICLK), .D(BIST_RDATA_T1160_4), .S(TRST_
        ), .Q(BIST_RDATA_T_4) );
    zdffqsb BIST_RDATA_reg_22 ( .CK(PCICLK), .D(BIST_RDATA1122_22), .S(TRST_), 
        .Q(BIST_RDATA_22) );
    zdffqsb BIST_WDATA_reg_26 ( .CK(PCICLK), .D(BIST_WDATA734_26), .S(TRST_), 
        .Q(BIST_WDATA_26) );
    zdffqsb BIST_RDATA_reg_6 ( .CK(PCICLK), .D(BIST_RDATA1122_6), .S(TRST_), 
        .Q(BIST_RDATA_6) );
    zdffqsb BIST_RDATA_T_reg_12 ( .CK(PCICLK), .D(BIST_RDATA_T1160_12), .S(
        TRST_), .Q(BIST_RDATA_T_12) );
    zdffqrb BIST_RDATA_T_reg_27 ( .CK(PCICLK), .D(BIST_RDATA_T1160_27), .R(
        TRST_), .Q(BIST_RDATA_T_27) );
    zdffqsb BIST_WDATA_reg_2 ( .CK(PCICLK), .D(BIST_WDATA734_2), .S(TRST_), 
        .Q(BIST_WDATA_2) );
    zdffqrb BIST_WDATA_reg_13 ( .CK(PCICLK), .D(BIST_WDATA734_13), .R(TRST_), 
        .Q(BIST_WDATA_13) );
    zdffqrb BIST_RDATA_reg_17 ( .CK(PCICLK), .D(BIST_RDATA1122_17), .R(TRST_), 
        .Q(BIST_RDATA_17) );
    zdffqsb BIST_RDATA_reg_30 ( .CK(PCICLK), .D(BIST_RDATA1122_30), .S(TRST_), 
        .Q(BIST_RDATA_30) );
    zdffqsb BIST_RDATA_reg_10 ( .CK(PCICLK), .D(BIST_RDATA1122_10), .S(TRST_), 
        .Q(BIST_RDATA_10) );
    zdffqsb BIST_WDATA_reg_28 ( .CK(PCICLK), .D(BIST_WDATA734_28), .S(TRST_), 
        .Q(BIST_WDATA_28) );
    zdffqsb BIST_RDATA_reg_8 ( .CK(PCICLK), .D(BIST_RDATA1122_8), .S(TRST_), 
        .Q(BIST_RDATA_8) );
    zdffqsb BIST_WDATA_reg_14 ( .CK(PCICLK), .D(BIST_WDATA734_14), .S(TRST_), 
        .Q(BIST_WDATA_14) );
    zdffqrb BIST_WDATA_reg_5 ( .CK(PCICLK), .D(BIST_WDATA734_5), .R(TRST_), 
        .Q(BIST_WDATA_5) );
    zdffqsb BIST_RDATA_T_reg_20 ( .CK(PCICLK), .D(BIST_RDATA_T1160_20), .S(
        TRST_), .Q(BIST_RDATA_T_20) );
    zdffqrb BIST_ERR_S_reg ( .CK(PCICLK), .D(BIST_ERR_S1235), .R(TRST_), .Q(
        BIST_ERR_S) );
    zdffqrb BIST_RDATA_reg_19 ( .CK(PCICLK), .D(BIST_RDATA1122_19), .R(TRST_), 
        .Q(BIST_RDATA_19) );
    zdffqrb BIST_RDATA_T_reg_15 ( .CK(PCICLK), .D(BIST_RDATA_T1160_15), .R(
        TRST_), .Q(BIST_RDATA_T_15) );
    zdffqrb BIST_WDATA_reg_21 ( .CK(PCICLK), .D(BIST_WDATA734_21), .R(TRST_), 
        .Q(BIST_WDATA_21) );
    zdffqrb BIST_RDATA_reg_1 ( .CK(PCICLK), .D(BIST_RDATA1122_1), .R(TRST_), 
        .Q(BIST_RDATA_1) );
    zdffqrb BIST_RDATA_T_reg_3 ( .CK(PCICLK), .D(BIST_RDATA_T1160_3), .R(TRST_
        ), .Q(BIST_RDATA_T_3) );
    zdffqrb BIST_RDATA_T_reg_29 ( .CK(PCICLK), .D(BIST_RDATA_T1160_29), .R(
        TRST_), .Q(BIST_RDATA_T_29) );
    zdffqrb BIST_RDATA_reg_25 ( .CK(PCICLK), .D(BIST_RDATA1122_25), .R(TRST_), 
        .Q(BIST_RDATA_25) );
    zdffqrb BIST_RDATA_T_reg_21 ( .CK(PCICLK), .D(BIST_RDATA_T1160_21), .R(
        TRST_), .Q(BIST_RDATA_T_21) );
    zdffqrb BIST_RUN_T_reg ( .CK(PCICLK), .D(BIST_RUN), .R(TRST_), .Q(
        BIST_RUN_T) );
    zdffqrb BIST_WDATA_reg_15 ( .CK(PCICLK), .D(BIST_WDATA734_15), .R(TRST_), 
        .Q(BIST_WDATA_15) );
    zdffqsb BIST_WDATA_reg_4 ( .CK(PCICLK), .D(BIST_WDATA734_4), .S(TRST_), 
        .Q(BIST_WDATA_4) );
    zdffqrb BIST_RUN_C_reg ( .CK(PCICLK), .D(BIST_RUN_C346), .R(TRST_), .Q(
        BIST_RUN_C) );
    zdffqrb BIST_WDATA_reg_29 ( .CK(PCICLK), .D(BIST_WDATA734_29), .R(TRST_), 
        .Q(BIST_WDATA_29) );
    zdffqrb BIST_RDATA_reg_9 ( .CK(PCICLK), .D(BIST_RDATA1122_9), .R(TRST_), 
        .Q(BIST_RDATA_9) );
    zdffqrb BIST_RDATA_reg_11 ( .CK(PCICLK), .D(BIST_RDATA1122_11), .R(TRST_), 
        .Q(BIST_RDATA_11) );
    zdffqsb BIST_RDATA_T_reg_2 ( .CK(PCICLK), .D(BIST_RDATA_T1160_2), .S(TRST_
        ), .Q(BIST_RDATA_T_2) );
    zdffqsb BIST_RDATA_T_reg_28 ( .CK(PCICLK), .D(BIST_RDATA_T1160_28), .S(
        TRST_), .Q(BIST_RDATA_T_28) );
    zdffqrb_ SRAM_R_T_reg ( .CK(PCICLK), .D(SRAM_R_T1481), .R(TRST_), .Q(
        SRAM_R_T) );
    zdffqsb BIST_RDATA_reg_24 ( .CK(PCICLK), .D(BIST_RDATA1122_24), .S(TRST_), 
        .Q(BIST_RDATA_24) );
    zdffqsb BIST_WDATA_reg_20 ( .CK(PCICLK), .D(BIST_WDATA734_20), .S(TRST_), 
        .Q(BIST_WDATA_20) );
    zdffqsb BIST_RDATA_reg_0 ( .CK(PCICLK), .D(BIST_RDATA1122_0), .S(TRST_), 
        .Q(BIST_RDATA_0) );
    zdffqsb BIST_RDATA_reg_18 ( .CK(PCICLK), .D(BIST_RDATA1122_18), .S(TRST_), 
        .Q(BIST_RDATA_18) );
    zdffqsb BIST_RDATA_T_reg_14 ( .CK(PCICLK), .D(BIST_RDATA_T1160_14), .S(
        TRST_), .Q(BIST_RDATA_T_14) );
    zdffqrb BIST_RDATA_T_reg_13 ( .CK(PCICLK), .D(BIST_RDATA_T1160_13), .R(
        TRST_), .Q(BIST_RDATA_T_13) );
    zdffqrb BIST_WDATA_reg_27 ( .CK(PCICLK), .D(BIST_WDATA734_27), .R(TRST_), 
        .Q(BIST_WDATA_27) );
    zdffqrb BIST_RDATA_reg_7 ( .CK(PCICLK), .D(BIST_RDATA1122_7), .R(TRST_), 
        .Q(BIST_RDATA_7) );
    zdffqrb BIST_RDATA_T_reg_5 ( .CK(PCICLK), .D(BIST_RDATA_T1160_5), .R(TRST_
        ), .Q(BIST_RDATA_T_5) );
    zdffqrb BIST_RDATA_reg_23 ( .CK(PCICLK), .D(BIST_RDATA1122_23), .R(TRST_), 
        .Q(BIST_RDATA_23) );
    zdffqsb BIST_RDATA_reg_16 ( .CK(PCICLK), .D(BIST_RDATA1122_16), .S(TRST_), 
        .Q(BIST_RDATA_16) );
    zdffqrb BIST_RDATA_reg_31 ( .CK(PCICLK), .D(BIST_RDATA1122_31), .R(TRST_), 
        .Q(BIST_RDATA_31) );
    zdffqsb BIST_WDATA_reg_12 ( .CK(PCICLK), .D(BIST_WDATA734_12), .S(TRST_), 
        .Q(BIST_WDATA_12) );
    zdffqrb BIST_WDATA_reg_3 ( .CK(PCICLK), .D(BIST_WDATA734_3), .R(TRST_), 
        .Q(BIST_WDATA_3) );
    zdffqsb BIST_RDATA_T_reg_26 ( .CK(PCICLK), .D(BIST_RDATA_T1160_26), .S(
        TRST_), .Q(BIST_RDATA_T_26) );
    zdffqrb_ DATARDY_reg ( .CK(PCICLK), .D(n2446), .R(TRST_), .Q(DATARDY) );
    zdffqrb BIST_RDATA_reg_21 ( .CK(PCICLK), .D(BIST_RDATA1122_21), .R(TRST_), 
        .Q(BIST_RDATA_21) );
    zdffqrb BIST_RDATA_T_reg_7 ( .CK(PCICLK), .D(BIST_RDATA_T1160_7), .R(TRST_
        ), .Q(BIST_RDATA_T_7) );
    zdffqrb BIST_WDATA_reg_19 ( .CK(PCICLK), .D(BIST_WDATA734_19), .R(TRST_), 
        .Q(BIST_WDATA_19) );
    zdffqsb BIST_WDATA_reg_8 ( .CK(PCICLK), .D(BIST_WDATA734_8), .S(TRST_), 
        .Q(BIST_WDATA_8) );
    zdffqrb BIST_RDATA_reg_5 ( .CK(PCICLK), .D(BIST_RDATA1122_5), .R(TRST_), 
        .Q(BIST_RDATA_5) );
    zdffqrb BIST_WDATA_reg_25 ( .CK(PCICLK), .D(BIST_WDATA734_25), .R(TRST_), 
        .Q(BIST_WDATA_25) );
    zdffqrb BIST_RDATA_T_reg_11 ( .CK(PCICLK), .D(BIST_RDATA_T1160_11), .R(
        TRST_), .Q(BIST_RDATA_T_11) );
    zdffqrb_ BIST_WR_reg ( .CK(PCICLK), .D(BIST_WR1405), .R(TRST_), .Q(BIST_WR
        ) );
    zdffqrb_ BIST_RD_T_reg ( .CK(PCICLK), .D(BIST_RD_T1359), .R(TRST_), .Q(
        BIST_RD_T) );
    zivb U1159 ( .A(BIST_RD_T), .Y(n2178) );
    zdffqsb BIST_RDATA_reg_28 ( .CK(PCICLK), .D(BIST_RDATA1122_28), .S(TRST_), 
        .Q(BIST_RDATA_28) );
    zdffqsb BIST_RDATA_T_reg_24 ( .CK(PCICLK), .D(BIST_RDATA_T1160_24), .S(
        TRST_), .Q(BIST_RDATA_T_24) );
    zdffqrb BIST_WDATA_reg_1 ( .CK(PCICLK), .D(BIST_WDATA734_1), .R(TRST_), 
        .Q(BIST_WDATA_1) );
    zdffqsb BIST_WDATA_reg_10 ( .CK(PCICLK), .D(BIST_WDATA734_10), .S(TRST_), 
        .Q(BIST_WDATA_10) );
    zdffqsb BIST_RDATA_T_reg_18 ( .CK(PCICLK), .D(BIST_RDATA_T1160_18), .S(
        TRST_), .Q(BIST_RDATA_T_18) );
    zdffqrb_ SRAM_W_T_reg ( .CK(PCICLK), .D(SRAM_W_T1443), .R(TRST_), .Q(
        SRAM_W_T) );
    zdffqsb BIST_RDATA_reg_14 ( .CK(PCICLK), .D(BIST_RDATA1122_14), .S(TRST_), 
        .Q(BIST_RDATA_14) );
    zdffqrb BIST_RDATA_reg_13 ( .CK(PCICLK), .D(BIST_RDATA1122_13), .R(TRST_), 
        .Q(BIST_RDATA_13) );
    zdffqsb BIST_WDATA_reg_30 ( .CK(PCICLK), .D(BIST_WDATA734_30), .S(TRST_), 
        .Q(BIST_WDATA_30) );
    zdffqrb BIST_WDATA_reg_17 ( .CK(PCICLK), .D(BIST_WDATA734_17), .R(TRST_), 
        .Q(BIST_WDATA_17) );
    zdffqsb BIST_WDATA_reg_6 ( .CK(PCICLK), .D(BIST_WDATA734_6), .S(TRST_), 
        .Q(BIST_WDATA_6) );
    zdffqrb BIST_RDATA_T_reg_9 ( .CK(PCICLK), .D(BIST_RDATA_T1160_9), .R(TRST_
        ), .Q(BIST_RDATA_T_9) );
    zdffqrb BIST_RDATA_T_reg_23 ( .CK(PCICLK), .D(BIST_RDATA_T1160_23), .R(
        TRST_), .Q(BIST_RDATA_T_23) );
    zdffqrb BIST_RDATA_T_reg_31 ( .CK(PCICLK), .D(BIST_RDATA_T1160_31), .R(
        TRST_), .Q(BIST_RDATA_T_31) );
    zdffqsb BIST_RDATA_T_reg_16 ( .CK(PCICLK), .D(BIST_RDATA_T1160_16), .S(
        TRST_), .Q(BIST_RDATA_T_16) );
    zdffqsb BIST_WDATA_reg_22 ( .CK(PCICLK), .D(BIST_WDATA734_22), .S(TRST_), 
        .Q(BIST_WDATA_22) );
    zdffqsb BIST_RDATA_reg_2 ( .CK(PCICLK), .D(BIST_RDATA1122_2), .S(TRST_), 
        .Q(BIST_RDATA_2) );
    zdffqsb BIST_RDATA_reg_26 ( .CK(PCICLK), .D(BIST_RDATA1122_26), .S(TRST_), 
        .Q(BIST_RDATA_26) );
    zdffqsb BIST_RDATA_T_reg_0 ( .CK(PCICLK), .D(BIST_RDATA_T1160_0), .S(TRST_
        ), .Q(BIST_RDATA_T_0) );
    zdffqsb BIST_RDATA_T_reg_8 ( .CK(PCICLK), .D(BIST_RDATA_T1160_8), .S(TRST_
        ), .Q(BIST_RDATA_T_8) );
    zdffqsb BIST_RDATA_T_reg_22 ( .CK(PCICLK), .D(BIST_RDATA_T1160_22), .S(
        TRST_), .Q(BIST_RDATA_T_22) );
    zdffqrb BIST_WDATA_reg_31 ( .CK(PCICLK), .D(BIST_WDATA734_31), .R(TRST_), 
        .Q(BIST_WDATA_31) );
    zdffqsb BIST_WDATA_reg_16 ( .CK(PCICLK), .D(BIST_WDATA734_16), .S(TRST_), 
        .Q(BIST_WDATA_16) );
    zdffqrb BIST_WDATA_reg_7 ( .CK(PCICLK), .D(BIST_WDATA734_7), .R(TRST_), 
        .Q(BIST_WDATA_7) );
    zdffqsb BIST_RDATA_reg_12 ( .CK(PCICLK), .D(BIST_RDATA1122_12), .S(TRST_), 
        .Q(BIST_RDATA_12) );
    zdffqrb BIST_RDATA_reg_27 ( .CK(PCICLK), .D(BIST_RDATA1122_27), .R(TRST_), 
        .Q(BIST_RDATA_27) );
    zdffqrb BIST_RDATA_T_reg_1 ( .CK(PCICLK), .D(BIST_RDATA_T1160_1), .R(TRST_
        ), .Q(BIST_RDATA_T_1) );
    zdffqrb BIST_RDATA_reg_3 ( .CK(PCICLK), .D(BIST_RDATA1122_3), .R(TRST_), 
        .Q(BIST_RDATA_3) );
    zdffqrb_ RPOP_reg ( .CK(PCICLK), .D(RPOP187), .R(TRST_), .Q(RPOP) );
    zdffqrb BIST_WDATA_reg_23 ( .CK(PCICLK), .D(BIST_WDATA734_23), .R(TRST_), 
        .Q(BIST_WDATA_23) );
    zdffqsb BIST_RDATA_T_reg_30 ( .CK(PCICLK), .D(BIST_RDATA_T1160_30), .S(
        TRST_), .Q(BIST_RDATA_T_30) );
    zdffqrb BIST_RDATA_T_reg_17 ( .CK(PCICLK), .D(BIST_RDATA_T1160_17), .R(
        TRST_), .Q(BIST_RDATA_T_17) );
    zdffrb_ BIST_RD_reg ( .CK(PCICLK), .D(BIST_RD1353), .R(TRST_), .Q(BIST_RD), 
        .QN(n2214) );
    zdffqsb BIST_RDATA_T_reg_10 ( .CK(PCICLK), .D(BIST_RDATA_T1160_10), .S(
        TRST_), .Q(BIST_RDATA_T_10) );
    zdffqsb BIST_WDATA_reg_24 ( .CK(PCICLK), .D(BIST_WDATA734_24), .S(TRST_), 
        .Q(BIST_WDATA_24) );
    zdffqsb BIST_RDATA_reg_4 ( .CK(PCICLK), .D(BIST_RDATA1122_4), .S(TRST_), 
        .Q(BIST_RDATA_4) );
    zdffqsb BIST_WDATA_reg_18 ( .CK(PCICLK), .D(BIST_WDATA734_18), .S(TRST_), 
        .Q(BIST_WDATA_18) );
    zdffqrb BIST_WDATA_reg_9 ( .CK(PCICLK), .D(BIST_WDATA734_9), .R(TRST_), 
        .Q(BIST_WDATA_9) );
    zdffqsb BIST_RDATA_reg_20 ( .CK(PCICLK), .D(BIST_RDATA1122_20), .S(TRST_), 
        .Q(BIST_RDATA_20) );
    zdffqsb BIST_RDATA_T_reg_6 ( .CK(PCICLK), .D(BIST_RDATA_T1160_6), .S(TRST_
        ), .Q(BIST_RDATA_T_6) );
    zdffqrb BIST_RDATA_T_reg_19 ( .CK(PCICLK), .D(BIST_RDATA_T1160_19), .R(
        TRST_), .Q(BIST_RDATA_T_19) );
    zdffqrb BIST_RDATA_reg_15 ( .CK(PCICLK), .D(BIST_RDATA1122_15), .R(TRST_), 
        .Q(BIST_RDATA_15) );
    zdffqrb BIST_CMP_reg ( .CK(PCICLK), .D(RD), .R(TRST_), .Q(BIST_CMP) );
    zdffqrb BIST_WDATA_reg_11 ( .CK(PCICLK), .D(BIST_WDATA734_11), .R(TRST_), 
        .Q(BIST_WDATA_11) );
    zdffqsb BIST_WDATA_reg_0 ( .CK(PCICLK), .D(BIST_WDATA734_0), .S(TRST_), 
        .Q(BIST_WDATA_0) );
    zdffqrb BIST_RDATA_reg_29 ( .CK(PCICLK), .D(BIST_RDATA1122_29), .R(TRST_), 
        .Q(BIST_RDATA_29) );
    zdffqrb BIST_RDATA_T_reg_25 ( .CK(PCICLK), .D(BIST_RDATA_T1160_25), .R(
        TRST_), .Q(BIST_RDATA_T_25) );
    znr2b U1160 ( .A(n2231), .B(n2248), .Y(n1950) );
    znr3b U1161 ( .A(n2225), .B(n2230), .C(n2269), .Y(n1951) );
    znr3b U1162 ( .A(n2223), .B(n2230), .C(n2270), .Y(n1952) );
    znr3b U1163 ( .A(BISTSM_4), .B(n2232), .C(n2221), .Y(n1953) );
    znr4b U1164 ( .A(n2225), .B(n2226), .C(BISTSM_6), .D(n2224), .Y(n1954) );
    znr3b U1165 ( .A(BISTSM_2), .B(n2222), .C(n2221), .Y(n1955) );
    znr4b U1166 ( .A(n2014), .B(n2228), .C(BISTSM_8), .D(n2016), .Y(n1956) );
    znr4b U1167 ( .A(n2225), .B(n2227), .C(BISTSM_3), .D(n2224), .Y(n1957) );
    znr2b U1168 ( .A(n2211), .B(n2212), .Y(n1958) );
    zaoi22b U1169 ( .A(n2376), .B(BIST_WADDR_7), .C(BIST_WADDRNXT440_7), .D(
        n2192), .Y(n1959) );
    znr3b U1170 ( .A(n2178), .B(n2377), .C(BIST_REMPTY), .Y(n1960) );
    zaoi22b U1171 ( .A(n2375), .B(BIST_RADDR_0), .C(BIST_RADDRNXT829_0), .D(
        n2199), .Y(n1961) );
    zaoi22b U1172 ( .A(n2375), .B(BIST_RADDR_7), .C(BIST_RADDRNXT829_7), .D(
        n2199), .Y(n1962) );
    zmux21hb U1173 ( .A(n2369), .B(BISTSMNXT_3), .S(n2378), .Y(n1963) );
    zmux21hb U1174 ( .A(n2369), .B(BISTSMNXT_3), .S(n1959), .Y(n1964) );
    zmux21hb U1175 ( .A(n2369), .B(BISTSMNXT_3), .S(n2379), .Y(n1965) );
    zmux21hb U1176 ( .A(n2369), .B(BISTSMNXT_3), .S(n2380), .Y(n1966) );
    zmux21hb U1177 ( .A(n2373), .B(n2381), .S(n2383), .Y(n1967) );
    zmux21hb U1178 ( .A(n2373), .B(n2381), .S(n1962), .Y(n1968) );
    zmux21hb U1179 ( .A(n2373), .B(n2381), .S(n2384), .Y(n1969) );
    zmux21hb U1180 ( .A(n2373), .B(n2381), .S(n2385), .Y(n1970) );
    zor2b U1181 ( .A(n2021), .B(n2022), .Y(_cell_830_U3_Z_0) );
    zivb U1182 ( .A(_cell_830_U3_Z_0), .Y(n2256) );
    zivb U1183 ( .A(n2235), .Y(_cell_830_U14_Z_0) );
    zao21b U1184 ( .A(BISTSMNXT_5), .B(n2236), .C(n2237), .Y(n2235) );
    ziv11d U1185 ( .A(BIST_RUN), .Y(n1971), .Z(n1972) );
    zivb U1186 ( .A(n2393), .Y(n2386) );
    zivb U1187 ( .A(n2393), .Y(n2387) );
    zivb U1188 ( .A(n2395), .Y(n2390) );
    zivb U1189 ( .A(n2394), .Y(n2388) );
    zivb U1190 ( .A(n2397), .Y(n2392) );
    zivb U1191 ( .A(n2396), .Y(n2391) );
    zivb U1192 ( .A(n2394), .Y(n2389) );
    zivb U1193 ( .A(n2288), .Y(n2393) );
    zivb U1194 ( .A(n2288), .Y(n2396) );
    zivb U1195 ( .A(n2288), .Y(n2397) );
    zivb U1196 ( .A(n2259), .Y(n2288) );
    zivb U1197 ( .A(n2288), .Y(n2394) );
    zivb U1198 ( .A(n2288), .Y(n2395) );
    zbfb U1199 ( .A(n2289), .Y(n2403) );
    zbfb U1200 ( .A(n2289), .Y(n2398) );
    zbfb U1201 ( .A(n2289), .Y(n2399) );
    zbfb U1202 ( .A(n2289), .Y(n2401) );
    zivb U1203 ( .A(n2286), .Y(n2289) );
    zbfb U1204 ( .A(n2289), .Y(n2402) );
    zbfb U1205 ( .A(n2289), .Y(n2400) );
    zor2d U1206 ( .A(n2178), .B(n2194), .Y(n2285) );
    zivb U1207 ( .A(n2407), .Y(n2405) );
    zivb U1208 ( .A(n2407), .Y(n2406) );
    zivb U1209 ( .A(n2407), .Y(n2404) );
    zivb U1210 ( .A(n2285), .Y(n2407) );
    zivb U1211 ( .A(n2283), .Y(n1973) );
    zao22b U1212 ( .A(n2284), .B(BISTSMNXT_4), .C(BISTSMNXT_6), .D(BIST_RD_T), 
        .Y(n2283) );
    zbfb U1213 ( .A(n1973), .Y(n2412) );
    zbfb U1214 ( .A(n1973), .Y(n2409) );
    zbfb U1215 ( .A(n1973), .Y(n2411) );
    zbfb U1216 ( .A(n1973), .Y(n2408) );
    zbfb U1217 ( .A(n1973), .Y(n2410) );
    zivb U1218 ( .A(n2423), .Y(n2414) );
    zivb U1219 ( .A(n2423), .Y(n2413) );
    zivb U1220 ( .A(n2425), .Y(n2417) );
    zivb U1221 ( .A(n2425), .Y(n2418) );
    zivb U1222 ( .A(n2427), .Y(n2422) );
    zivb U1223 ( .A(n2427), .Y(n2421) );
    zivb U1224 ( .A(n2426), .Y(n2419) );
    zivb U1225 ( .A(n2426), .Y(n2420) );
    zivb U1226 ( .A(n2424), .Y(n2415) );
    zivb U1227 ( .A(n2424), .Y(n2416) );
    zivb U1228 ( .A(n2275), .Y(n2423) );
    zivb U1229 ( .A(n2275), .Y(n2425) );
    zivb U1230 ( .A(n2275), .Y(n2427) );
    zivb U1231 ( .A(n2240), .Y(n2275) );
    zivb U1232 ( .A(n2275), .Y(n2424) );
    zivb U1233 ( .A(n2275), .Y(n2426) );
    zivb U1234 ( .A(n2433), .Y(n2432) );
    zivb U1235 ( .A(n2433), .Y(n2429) );
    zivb U1236 ( .A(n2433), .Y(n2431) );
    zivb U1237 ( .A(n2433), .Y(n2428) );
    zivb U1238 ( .A(n2433), .Y(n2430) );
    zcx3b U1239 ( .A(n2179), .B(BISTSM_1), .C(n2371), .D(n2372), .Y(n2276) );
    zivb U1240 ( .A(n2276), .Y(n2433) );
    zbfb U1241 ( .A(n2274), .Y(n2435) );
    zbfb U1242 ( .A(n2274), .Y(n2438) );
    zbfb U1243 ( .A(n2274), .Y(n2434) );
    zivb U1244 ( .A(n2273), .Y(n2274) );
    zbfb U1245 ( .A(n2274), .Y(n2439) );
    zbfb U1246 ( .A(n2274), .Y(n2436) );
    zbfb U1247 ( .A(n2274), .Y(n2437) );
    zivb U1248 ( .A(n2272), .Y(n1974) );
    zao22b U1249 ( .A(BISTSMNXT_6), .B(n2179), .C(BISTSMNXT_4), .D(n2236), .Y(
        n2272) );
    zbfb U1250 ( .A(n1974), .Y(n2444) );
    zbfb U1251 ( .A(n1974), .Y(n2441) );
    zbfb U1252 ( .A(n1974), .Y(n2443) );
    zbfb U1253 ( .A(n1974), .Y(n2440) );
    zbfb U1254 ( .A(n1974), .Y(n2442) );
    zivc U1255 ( .A(n1977), .Y(n1978) );
    zan3b U1256 ( .A(SRAM_RUN), .B(n2213), .C(n1958), .Y(n1975) );
    zivc U1257 ( .A(n1971), .Y(n1976) );
    zivb U1258 ( .A(n1971), .Y(n1736) );
    zivb U1259 ( .A(n1975), .Y(n1977) );
    zivb U1260 ( .A(n1977), .Y(n1979) );
    zivb U1261 ( .A(n2213), .Y(n1980) );
    zivb U1262 ( .A(SRAM_RUN_T), .Y(n2213) );
    zdffqrb SRAM_RUN_T_reg ( .CK(PCICLK), .D(n1978), .R(TRST_), .Q(SRAM_RUN_T)
         );
    zdffqd RADDR_ATPG_reg_8 ( .CK(ATPG_CLK), .D(RADDR[8]), .Q(RADDR_ATPG[8])
         );
    zdffqd RADDR_ATPG_reg_7 ( .CK(ATPG_CLK), .D(RADDR[7]), .Q(RADDR_ATPG[7])
         );
    zdffqd RADDR_ATPG_reg_6 ( .CK(ATPG_CLK), .D(RADDR[6]), .Q(RADDR_ATPG[6])
         );
    zdffqd RADDR_ATPG_reg_5 ( .CK(ATPG_CLK), .D(RADDR[5]), .Q(RADDR_ATPG[5])
         );
    zdffqd RADDR_ATPG_reg_4 ( .CK(ATPG_CLK), .D(RADDR[4]), .Q(RADDR_ATPG[4])
         );
    zdffqd RADDR_ATPG_reg_3 ( .CK(ATPG_CLK), .D(RADDR[3]), .Q(RADDR_ATPG[3])
         );
    zdffqd RADDR_ATPG_reg_2 ( .CK(ATPG_CLK), .D(RADDR[2]), .Q(RADDR_ATPG[2])
         );
    zdffqd RADDR_ATPG_reg_1 ( .CK(ATPG_CLK), .D(RADDR[1]), .Q(RADDR_ATPG[1])
         );
    zdffqd RADDR_ATPG_reg_0 ( .CK(ATPG_CLK), .D(RADDR[0]), .Q(RADDR_ATPG[0])
         );
    zdffqd WADDR_ATPG_reg_8 ( .CK(ATPG_CLK), .D(WADDR[8]), .Q(WADDR_ATPG[8])
         );
    zdffqd WADDR_ATPG_reg_7 ( .CK(ATPG_CLK), .D(WADDR[7]), .Q(WADDR_ATPG[7])
         );
    zdffqd WADDR_ATPG_reg_6 ( .CK(ATPG_CLK), .D(WADDR[6]), .Q(WADDR_ATPG[6])
         );
    zdffqd WADDR_ATPG_reg_5 ( .CK(ATPG_CLK), .D(WADDR[5]), .Q(WADDR_ATPG[5])
         );
    zdffqd WADDR_ATPG_reg_4 ( .CK(ATPG_CLK), .D(WADDR[4]), .Q(WADDR_ATPG[4])
         );
    zdffqd WADDR_ATPG_reg_3 ( .CK(ATPG_CLK), .D(WADDR[3]), .Q(WADDR_ATPG[3])
         );
    zdffqd WADDR_ATPG_reg_2 ( .CK(ATPG_CLK), .D(WADDR[2]), .Q(WADDR_ATPG[2])
         );
    zdffqd WADDR_ATPG_reg_1 ( .CK(ATPG_CLK), .D(WADDR[1]), .Q(WADDR_ATPG[1])
         );
    zdffqd WADDR_ATPG_reg_0 ( .CK(ATPG_CLK), .D(WADDR_ATPG1549_0), .Q(
        WADDR_ATPG[0]) );
    zdffqd MDI_ATPG_reg_31 ( .CK(ATPG_CLK), .D(MDI[31]), .Q(MDI_ATPG[31]) );
    zdffqd MDI_ATPG_reg_30 ( .CK(ATPG_CLK), .D(MDI[30]), .Q(MDI_ATPG[30]) );
    zdffqd MDI_ATPG_reg_29 ( .CK(ATPG_CLK), .D(MDI[29]), .Q(MDI_ATPG[29]) );
    zdffqd MDI_ATPG_reg_28 ( .CK(ATPG_CLK), .D(MDI[28]), .Q(MDI_ATPG[28]) );
    zdffqd MDI_ATPG_reg_27 ( .CK(ATPG_CLK), .D(MDI[27]), .Q(MDI_ATPG[27]) );
    zdffqd MDI_ATPG_reg_26 ( .CK(ATPG_CLK), .D(MDI[26]), .Q(MDI_ATPG[26]) );
    zdffqd MDI_ATPG_reg_25 ( .CK(ATPG_CLK), .D(MDI[25]), .Q(MDI_ATPG[25]) );
    zdffqd MDI_ATPG_reg_24 ( .CK(ATPG_CLK), .D(MDI[24]), .Q(MDI_ATPG[24]) );
    zdffqd MDI_ATPG_reg_23 ( .CK(ATPG_CLK), .D(MDI[23]), .Q(MDI_ATPG[23]) );
    zdffqd MDI_ATPG_reg_22 ( .CK(ATPG_CLK), .D(MDI[22]), .Q(MDI_ATPG[22]) );
    zdffqd MDI_ATPG_reg_21 ( .CK(ATPG_CLK), .D(MDI[21]), .Q(MDI_ATPG[21]) );
    zdffqd MDI_ATPG_reg_20 ( .CK(ATPG_CLK), .D(MDI[20]), .Q(MDI_ATPG[20]) );
    zdffqd MDI_ATPG_reg_19 ( .CK(ATPG_CLK), .D(MDI[19]), .Q(MDI_ATPG[19]) );
    zdffqd MDI_ATPG_reg_18 ( .CK(ATPG_CLK), .D(MDI[18]), .Q(MDI_ATPG[18]) );
    zdffqd MDI_ATPG_reg_17 ( .CK(ATPG_CLK), .D(MDI[17]), .Q(MDI_ATPG[17]) );
    zdffqd MDI_ATPG_reg_16 ( .CK(ATPG_CLK), .D(MDI[16]), .Q(MDI_ATPG[16]) );
    zdffqd MDI_ATPG_reg_15 ( .CK(ATPG_CLK), .D(MDI[15]), .Q(MDI_ATPG[15]) );
    zdffqd MDI_ATPG_reg_14 ( .CK(ATPG_CLK), .D(MDI[14]), .Q(MDI_ATPG[14]) );
    zdffqd MDI_ATPG_reg_13 ( .CK(ATPG_CLK), .D(MDI[13]), .Q(MDI_ATPG[13]) );
    zdffqd MDI_ATPG_reg_12 ( .CK(ATPG_CLK), .D(MDI[12]), .Q(MDI_ATPG[12]) );
    zdffqd MDI_ATPG_reg_11 ( .CK(ATPG_CLK), .D(MDI[11]), .Q(MDI_ATPG[11]) );
    zdffqd MDI_ATPG_reg_10 ( .CK(ATPG_CLK), .D(MDI[10]), .Q(MDI_ATPG[10]) );
    zdffqd MDI_ATPG_reg_9 ( .CK(ATPG_CLK), .D(MDI[9]), .Q(MDI_ATPG[9]) );
    zdffqd MDI_ATPG_reg_8 ( .CK(ATPG_CLK), .D(MDI[8]), .Q(MDI_ATPG[8]) );
    zdffqd MDI_ATPG_reg_7 ( .CK(ATPG_CLK), .D(MDI[7]), .Q(MDI_ATPG[7]) );
    zdffqd MDI_ATPG_reg_6 ( .CK(ATPG_CLK), .D(MDI[6]), .Q(MDI_ATPG[6]) );
    zdffqd MDI_ATPG_reg_5 ( .CK(ATPG_CLK), .D(MDI[5]), .Q(MDI_ATPG[5]) );
    zdffqd MDI_ATPG_reg_4 ( .CK(ATPG_CLK), .D(MDI[4]), .Q(MDI_ATPG[4]) );
    zdffqd MDI_ATPG_reg_3 ( .CK(ATPG_CLK), .D(MDI[3]), .Q(MDI_ATPG[3]) );
    zdffqd MDI_ATPG_reg_2 ( .CK(ATPG_CLK), .D(MDI[2]), .Q(MDI_ATPG[2]) );
    zdffqd MDI_ATPG_reg_1 ( .CK(ATPG_CLK), .D(MDI[1]), .Q(MDI_ATPG[1]) );
    zdffqd MDI_ATPG_reg_0 ( .CK(ATPG_CLK), .D(MDI[0]), .Q(MDI_ATPG[0]) );
    zfa1b r133_U1_5 ( .A(BIST_WADDR_5), .B(_cell_830_U14_Z_0), .CI(
        r133_carry_5), .CO(r133_carry_6), .S(BIST_WADDRNXT440_5) );
    zfa1b r133_U1_4 ( .A(BIST_WADDR_4), .B(_cell_830_U14_Z_0), .CI(
        r133_carry_4), .CO(r133_carry_5), .S(BIST_WADDRNXT440_4) );
    zfa1b r133_U1_3 ( .A(BIST_WADDR_3), .B(_cell_830_U14_Z_0), .CI(
        r133_carry_3), .CO(r133_carry_4), .S(BIST_WADDRNXT440_3) );
    zfa1b r133_U1_2 ( .A(BIST_WADDR_2), .B(_cell_830_U14_Z_0), .CI(
        r133_carry_2), .CO(r133_carry_3), .S(BIST_WADDRNXT440_2) );
    zfa1b r133_U1_7 ( .A(BIST_WADDR_7), .B(_cell_830_U14_Z_0), .CI(
        r133_carry_7), .CO(r133_carry_8), .S(BIST_WADDRNXT440_7) );
    zfa1b r133_U1_0 ( .A(BIST_WADDR_0), .B(_cell_830_U14_Z_0), .CI(n2235), 
        .CO(r133_carry_1), .S(BIST_WADDRNXT440_0) );
    zfa1b r133_U1_6 ( .A(BIST_WADDR_6), .B(_cell_830_U14_Z_0), .CI(
        r133_carry_6), .CO(r133_carry_7), .S(BIST_WADDRNXT440_6) );
    zfa1b r133_U1_1 ( .A(BIST_WADDR_1), .B(_cell_830_U14_Z_0), .CI(
        r133_carry_1), .CO(r133_carry_2), .S(BIST_WADDRNXT440_1) );
    zfa1b r143_U1_5 ( .A(BIST_RADDR_5), .B(_cell_830_U3_Z_0), .CI(r143_carry_5
        ), .CO(r143_carry_6), .S(BIST_RADDRNXT829_5) );
    zfa1b r143_U1_4 ( .A(BIST_RADDR_4), .B(_cell_830_U3_Z_0), .CI(r143_carry_4
        ), .CO(r143_carry_5), .S(BIST_RADDRNXT829_4) );
    zfa1b r143_U1_3 ( .A(BIST_RADDR_3), .B(_cell_830_U3_Z_0), .CI(r143_carry_3
        ), .CO(r143_carry_4), .S(BIST_RADDRNXT829_3) );
    zfa1b r143_U1_2 ( .A(BIST_RADDR_2), .B(_cell_830_U3_Z_0), .CI(r143_carry_2
        ), .CO(r143_carry_3), .S(BIST_RADDRNXT829_2) );
    zfa1b r143_U1_7 ( .A(BIST_RADDR_7), .B(_cell_830_U3_Z_0), .CI(r143_carry_7
        ), .CO(r143_carry_8), .S(BIST_RADDRNXT829_7) );
    zfa1b r143_U1_0 ( .A(BIST_RADDR_0), .B(_cell_830_U3_Z_0), .CI(n2256), .CO(
        r143_carry_1), .S(BIST_RADDRNXT829_0) );
    zfa1b r143_U1_6 ( .A(BIST_RADDR_6), .B(_cell_830_U3_Z_0), .CI(r143_carry_6
        ), .CO(r143_carry_7), .S(BIST_RADDRNXT829_6) );
    zfa1b r143_U1_1 ( .A(BIST_RADDR_1), .B(_cell_830_U3_Z_0), .CI(r143_carry_1
        ), .CO(r143_carry_2), .S(BIST_RADDRNXT829_1) );
    zinr2b U1263 ( .A(RMA[8]), .B(SLAVEMODE), .Y(n1983) );
    zao211b U1264 ( .A(BIST_WR), .B(n1736), .C(SRAM_W_T), .D(n2008), .Y(WR) );
    zan4b U1265 ( .A(BIST_CMP), .B(BIST_RUN_T), .C(n1740), .D(n2018), .Y(
        BIST_ERR_S1235) );
    zor3b U1266 ( .A(n2023), .B(n2024), .C(n2025), .Y(BIST_WDATA734_0) );
    zor3b U1267 ( .A(n2026), .B(n2027), .C(n1963), .Y(BIST_WDATA734_1) );
    zor3b U1268 ( .A(n2028), .B(n2029), .C(n2030), .Y(BIST_WDATA734_2) );
    zor3b U1269 ( .A(n2031), .B(n2032), .C(n1966), .Y(BIST_WDATA734_3) );
    zor3b U1270 ( .A(n2033), .B(n2034), .C(n2035), .Y(BIST_WDATA734_4) );
    zor3b U1271 ( .A(n2036), .B(n2037), .C(n1965), .Y(BIST_WDATA734_5) );
    zor3b U1272 ( .A(n2038), .B(n2039), .C(n2040), .Y(BIST_WDATA734_6) );
    zor3b U1273 ( .A(n2041), .B(n2042), .C(n1964), .Y(BIST_WDATA734_7) );
    zor3b U1274 ( .A(n2043), .B(n2044), .C(n2025), .Y(BIST_WDATA734_8) );
    zor3b U1275 ( .A(n2045), .B(n2046), .C(n1963), .Y(BIST_WDATA734_9) );
    zor3b U1276 ( .A(n2047), .B(n2048), .C(n2030), .Y(BIST_WDATA734_10) );
    zor3b U1277 ( .A(n2049), .B(n2050), .C(n1966), .Y(BIST_WDATA734_11) );
    zor3b U1278 ( .A(n2051), .B(n2052), .C(n2035), .Y(BIST_WDATA734_12) );
    zor3b U1279 ( .A(n2053), .B(n2054), .C(n1965), .Y(BIST_WDATA734_13) );
    zor3b U1280 ( .A(n2055), .B(n2056), .C(n2040), .Y(BIST_WDATA734_14) );
    zor3b U1281 ( .A(n2057), .B(n2058), .C(n1964), .Y(BIST_WDATA734_15) );
    zor3b U1282 ( .A(n2059), .B(n2060), .C(n2025), .Y(BIST_WDATA734_16) );
    zor3b U1283 ( .A(n2061), .B(n2062), .C(n1963), .Y(BIST_WDATA734_17) );
    zor3b U1284 ( .A(n2063), .B(n2064), .C(n2030), .Y(BIST_WDATA734_18) );
    zor3b U1285 ( .A(n2065), .B(n2066), .C(n1966), .Y(BIST_WDATA734_19) );
    zor3b U1286 ( .A(n2067), .B(n2068), .C(n2035), .Y(BIST_WDATA734_20) );
    zor3b U1287 ( .A(n2069), .B(n2070), .C(n1965), .Y(BIST_WDATA734_21) );
    zor3b U1288 ( .A(n2071), .B(n2072), .C(n2040), .Y(BIST_WDATA734_22) );
    zor3b U1289 ( .A(n2073), .B(n2074), .C(n1964), .Y(BIST_WDATA734_23) );
    zor3b U1290 ( .A(n2075), .B(n2076), .C(n2025), .Y(BIST_WDATA734_24) );
    zor3b U1291 ( .A(n2077), .B(n2078), .C(n1963), .Y(BIST_WDATA734_25) );
    zor3b U1292 ( .A(n2079), .B(n2080), .C(n2030), .Y(BIST_WDATA734_26) );
    zor3b U1293 ( .A(n2081), .B(n2082), .C(n1966), .Y(BIST_WDATA734_27) );
    zor3b U1294 ( .A(n2083), .B(n2084), .C(n2035), .Y(BIST_WDATA734_28) );
    zor3b U1295 ( .A(n2085), .B(n2086), .C(n1965), .Y(BIST_WDATA734_29) );
    zor3b U1296 ( .A(n2087), .B(n2088), .C(n2040), .Y(BIST_WDATA734_30) );
    zor3b U1297 ( .A(n2089), .B(n2090), .C(n1964), .Y(BIST_WDATA734_31) );
    zor3b U1298 ( .A(n2091), .B(n2092), .C(n2093), .Y(BIST_RDATA1122_0) );
    zor3b U1299 ( .A(n1967), .B(n2094), .C(n2095), .Y(BIST_RDATA1122_1) );
    zor3b U1300 ( .A(n2096), .B(n2097), .C(n2098), .Y(BIST_RDATA1122_2) );
    zor3b U1301 ( .A(n2099), .B(n2100), .C(n1970), .Y(BIST_RDATA1122_3) );
    zor3b U1302 ( .A(n2101), .B(n2102), .C(n2103), .Y(BIST_RDATA1122_4) );
    zor3b U1303 ( .A(n2104), .B(n2105), .C(n1969), .Y(BIST_RDATA1122_5) );
    zor3b U1304 ( .A(n2106), .B(n2107), .C(n2108), .Y(BIST_RDATA1122_6) );
    zor3b U1305 ( .A(n2109), .B(n2110), .C(n1968), .Y(BIST_RDATA1122_7) );
    zor3b U1306 ( .A(n2111), .B(n2112), .C(n2093), .Y(BIST_RDATA1122_8) );
    zor3b U1307 ( .A(n1967), .B(n2113), .C(n2114), .Y(BIST_RDATA1122_9) );
    zor3b U1308 ( .A(n2115), .B(n2116), .C(n2098), .Y(BIST_RDATA1122_10) );
    zor3b U1309 ( .A(n2117), .B(n2118), .C(n1970), .Y(BIST_RDATA1122_11) );
    zor3b U1310 ( .A(n2119), .B(n2120), .C(n2103), .Y(BIST_RDATA1122_12) );
    zor3b U1311 ( .A(n2121), .B(n2122), .C(n1969), .Y(BIST_RDATA1122_13) );
    zor3b U1312 ( .A(n2123), .B(n2124), .C(n2108), .Y(BIST_RDATA1122_14) );
    zor3b U1313 ( .A(n2125), .B(n2126), .C(n1968), .Y(BIST_RDATA1122_15) );
    zor3b U1314 ( .A(n2127), .B(n2128), .C(n2093), .Y(BIST_RDATA1122_16) );
    zor3b U1315 ( .A(n1967), .B(n2129), .C(n2130), .Y(BIST_RDATA1122_17) );
    zor3b U1316 ( .A(n2131), .B(n2132), .C(n2098), .Y(BIST_RDATA1122_18) );
    zor3b U1317 ( .A(n2133), .B(n2134), .C(n1970), .Y(BIST_RDATA1122_19) );
    zor3b U1318 ( .A(n2135), .B(n2136), .C(n2103), .Y(BIST_RDATA1122_20) );
    zor3b U1319 ( .A(n2137), .B(n2138), .C(n1969), .Y(BIST_RDATA1122_21) );
    zor3b U1320 ( .A(n2139), .B(n2140), .C(n2108), .Y(BIST_RDATA1122_22) );
    zor3b U1321 ( .A(n2141), .B(n2142), .C(n1968), .Y(BIST_RDATA1122_23) );
    zor3b U1322 ( .A(n2143), .B(n2144), .C(n2093), .Y(BIST_RDATA1122_24) );
    zor3b U1323 ( .A(n1967), .B(n2145), .C(n2146), .Y(BIST_RDATA1122_25) );
    zor3b U1324 ( .A(n2147), .B(n2148), .C(n2098), .Y(BIST_RDATA1122_26) );
    zor3b U1325 ( .A(n2149), .B(n2150), .C(n1970), .Y(BIST_RDATA1122_27) );
    zor3b U1326 ( .A(n2151), .B(n2152), .C(n2103), .Y(BIST_RDATA1122_28) );
    zor3b U1327 ( .A(n2153), .B(n2154), .C(n1969), .Y(BIST_RDATA1122_29) );
    zor3b U1328 ( .A(n2155), .B(n2156), .C(n2108), .Y(BIST_RDATA1122_30) );
    zor3b U1329 ( .A(n2157), .B(n2158), .C(n1968), .Y(BIST_RDATA1122_31) );
    zoai22d U1330 ( .A(ASYNCFIFO), .B(n2159), .C(n2160), .D(n2161), .Y(
        BIST_RADDR1065_8) );
    zoai22d U1331 ( .A(n2162), .B(n2159), .C(n1962), .D(n2161), .Y(
        BIST_RADDR1065_7) );
    zoai22d U1332 ( .A(ASYNCFIFO), .B(n2159), .C(n2170), .D(n2161), .Y(
        BIST_WADDR677_8) );
    zoai22d U1333 ( .A(n2162), .B(n2159), .C(n1959), .D(n2161), .Y(
        BIST_WADDR677_7) );
    zor6b U1334 ( .A(n2180), .B(n2181), .C(n2182), .D(n2183), .E(n2184), .F(
        n2185), .Y(n2179) );
    zinr2b U1335 ( .A(FPUSH), .B(SLAVE_ACT), .Y(n2008) );
    zoa21d U1336 ( .A(BISTSMNXT_3), .B(BISTSMNXT_6), .C(BIST_WUNDER), .Y(n2188
        ) );
    zor3b U1337 ( .A(BISTSMNXT_3), .B(n1952), .C(n2191), .Y(n2190) );
    zoa21d U1338 ( .A(BISTSM_6), .B(BISTSM_5), .C(n2009), .Y(n2197) );
    zoa21d U1339 ( .A(n2178), .B(BIST_RFULL), .C(BISTSMNXT_5), .Y(n2209) );
    zoa21d U1340 ( .A(n2178), .B(BIST_REMPTY), .C(n2191), .Y(n2210) );
    zor3b U1341 ( .A(BISTSM_2), .B(BISTSM_4), .C(BISTSM_0), .Y(n2016) );
    zor6b U1342 ( .A(BIST_RADDR_3), .B(BIST_RADDR_2), .C(BIST_RADDR_1), .D(
        BIST_RADDR_6), .E(BIST_RADDR_5), .F(BIST_RADDR_4), .Y(n2219) );
    zor4b U1343 ( .A(BISTSM_1), .B(BISTSM_3), .C(BISTSM_7), .D(BISTSM_6), .Y(
        n2014) );
    zor4b U1344 ( .A(BISTSM_5), .B(BISTSM_0), .C(BISTSM_8), .D(n2014), .Y(
        n2221) );
    zor4b U1345 ( .A(BIST_RADDR_7), .B(BIST_RADDR_8), .C(BIST_RADDR_0), .D(
        n2219), .Y(n2011) );
    zor3b U1346 ( .A(n2219), .B(n2220), .C(n2229), .Y(n2009) );
    zor5b U1347 ( .A(BISTSM_4), .B(BISTSM_2), .C(BISTSM_5), .D(BISTSM_3), .E(
        BISTSM_6), .Y(n2230) );
    zor3b U1348 ( .A(BISTSM_0), .B(BISTSM_1), .C(n2230), .Y(n2231) );
    zor3b U1349 ( .A(n1950), .B(n1951), .C(n1952), .Y(n2239) );
    zor5b U1350 ( .A(n1950), .B(n1951), .C(n2189), .D(BISTSMNXT_5), .E(n2190), 
        .Y(n2020) );
    zao211b U1351 ( .A(BISTSMNXT_5), .B(n2228), .C(n2247), .D(n2019), .Y(n2161
        ) );
    zoai22d U1352 ( .A(n2214), .B(n2258), .C(n2234), .D(n2022), .Y(n2259) );
    zao211b U1353 ( .A(BIST_RD), .B(n1976), .C(FPOP), .D(SRAM_R_T), .Y(n2265)
         );
    zor3b U1354 ( .A(n2209), .B(n2210), .C(n2287), .Y(n2286) );
    zor4b U1355 ( .A(n2217), .B(n2218), .C(n2215), .D(n2216), .Y(n2185) );
    zan4b U1356 ( .A(BISTSM_1), .B(n2234), .C(n2295), .D(n2296), .Y(n2010) );
    zor4b U1357 ( .A(n2253), .B(n2254), .C(n2251), .D(n2252), .Y(n2297) );
    zao222b U1358 ( .A(n2257), .B(n2189), .C(BISTSMNXT_3), .D(n2178), .E(n2298
        ), .F(n2239), .Y(n2287) );
    zor4b U1359 ( .A(n2317), .B(n2326), .C(n2299), .D(n2308), .Y(n2018) );
    zor3b U1360 ( .A(BIST_WFULL), .B(n2367), .C(n2368), .Y(n2277) );
    zoai22d U1361 ( .A(BIST_WUNDER), .B(n2377), .C(BIST_WFULL), .D(n2021), .Y(
        n2012) );
    zor6b U1362 ( .A(n2249), .B(n2250), .C(n2203), .D(n2220), .E(n2200), .F(
        n2297), .Y(n2015) );
    zor4b U1363 ( .A(BISTSM_1), .B(BISTSM_3), .C(n2198), .D(n2197), .Y(n2017)
         );
    zor3b U1364 ( .A(n2239), .B(n2189), .C(n2188), .Y(n2372) );
    zivb U1365 ( .A(RPOP), .Y(n2445) );
    zivb U1366 ( .A(n2445), .Y(n2446) );
endmodule


module FIFO_ATPG_MUX ( ATPG_ENI, DOUT, MDI_ATPG, MDO );
input  [31:0] DOUT;
output [31:0] MDO;
input  [31:0] MDI_ATPG;
input  ATPG_ENI;
    zymx24hb U12 ( .A1(DOUT[3]), .A2(DOUT[2]), .A3(DOUT[1]), .A4(DOUT[0]), 
        .B1(MDI_ATPG[3]), .B2(MDI_ATPG[2]), .B3(MDI_ATPG[1]), .B4(MDI_ATPG[0]), 
        .S(ATPG_ENI), .Y1(MDO[3]), .Y2(MDO[2]), .Y3(MDO[1]), .Y4(MDO[0]) );
    zymx24hb U13 ( .A1(DOUT[7]), .A2(DOUT[6]), .A3(DOUT[5]), .A4(DOUT[4]), 
        .B1(MDI_ATPG[7]), .B2(MDI_ATPG[6]), .B3(MDI_ATPG[5]), .B4(MDI_ATPG[4]), 
        .S(ATPG_ENI), .Y1(MDO[7]), .Y2(MDO[6]), .Y3(MDO[5]), .Y4(MDO[4]) );
    zymx24hb U14 ( .A1(DOUT[11]), .A2(DOUT[10]), .A3(DOUT[9]), .A4(DOUT[8]), 
        .B1(MDI_ATPG[11]), .B2(MDI_ATPG[10]), .B3(MDI_ATPG[9]), .B4(MDI_ATPG
        [8]), .S(ATPG_ENI), .Y1(MDO[11]), .Y2(MDO[10]), .Y3(MDO[9]), .Y4(MDO
        [8]) );
    zymx24hb U15 ( .A1(DOUT[15]), .A2(DOUT[14]), .A3(DOUT[13]), .A4(DOUT[12]), 
        .B1(MDI_ATPG[15]), .B2(MDI_ATPG[14]), .B3(MDI_ATPG[13]), .B4(MDI_ATPG
        [12]), .S(ATPG_ENI), .Y1(MDO[15]), .Y2(MDO[14]), .Y3(MDO[13]), .Y4(MDO
        [12]) );
    zymx24hb U16 ( .A1(DOUT[19]), .A2(DOUT[18]), .A3(DOUT[17]), .A4(DOUT[16]), 
        .B1(MDI_ATPG[19]), .B2(MDI_ATPG[18]), .B3(MDI_ATPG[17]), .B4(MDI_ATPG
        [16]), .S(ATPG_ENI), .Y1(MDO[19]), .Y2(MDO[18]), .Y3(MDO[17]), .Y4(MDO
        [16]) );
    zymx24hb U17 ( .A1(DOUT[23]), .A2(DOUT[22]), .A3(DOUT[21]), .A4(DOUT[20]), 
        .B1(MDI_ATPG[23]), .B2(MDI_ATPG[22]), .B3(MDI_ATPG[21]), .B4(MDI_ATPG
        [20]), .S(ATPG_ENI), .Y1(MDO[23]), .Y2(MDO[22]), .Y3(MDO[21]), .Y4(MDO
        [20]) );
    zymx24hb U18 ( .A1(DOUT[27]), .A2(DOUT[26]), .A3(DOUT[25]), .A4(DOUT[24]), 
        .B1(MDI_ATPG[27]), .B2(MDI_ATPG[26]), .B3(MDI_ATPG[25]), .B4(MDI_ATPG
        [24]), .S(ATPG_ENI), .Y1(MDO[27]), .Y2(MDO[26]), .Y3(MDO[25]), .Y4(MDO
        [24]) );
    zymx24hb U19 ( .A1(DOUT[31]), .A2(DOUT[30]), .A3(DOUT[29]), .A4(DOUT[28]), 
        .B1(MDI_ATPG[31]), .B2(MDI_ATPG[30]), .B3(MDI_ATPG[29]), .B4(MDI_ATPG
        [28]), .S(ATPG_ENI), .Y1(MDO[31]), .Y2(MDO[30]), .Y3(MDO[29]), .Y4(MDO
        [28]) );
endmodule


module DBG_FFCTL ( SRAM8_WE, DI, BUF_WE, BUF_DI, BUF_DAT1, BUF_DAT2, DBG_GO, 
    LATCHDAT, USBPOP, USBDAT, HOSTDAT, CLK60M, HRST_ );
input  [7:0] SRAM8_WE;
input  [31:0] DI;
output [7:0] BUF_WE;
output [31:0] BUF_DI;
input  [31:0] BUF_DAT2;
output [7:0] HOSTDAT;
input  [31:0] BUF_DAT1;
input  [7:0] USBDAT;
input  DBG_GO, LATCHDAT, USBPOP, CLK60M, HRST_;
    wire DBG_GO_T, SRAM8_WE_CLK60M177_6, SRAM8_WE_CLK60M_1, SPAREO6, 
        BUF_SEL139_2, BUF_SEL_2, SPAREO0_, BUF_SEL_5, BUF_SEL139_5, 
        SRAM8_WE_CLK60M_6, SPAREO1, BUF_SEL_4, SRAM8_WE_CLK60M177_1, 
        BUF_SEL139_4, SPAREO9, SRAM8_WE_CLK60M177_0, SRAM8_WE_CLK60M_7, 
        SPAREO0, SPAREO7, SRAM8_WE_CLK60M_0, SRAM8_WE_CLK60M177_7, BUF_SEL_3, 
        BUF_SEL139_3, SRAM8_WE_CLK60M177_5, SRAM8_WE_CLK60M_2, SPAREO5, 
        BUF_SEL_1, BUF_SEL139_1, BUF_SEL2_0, BUF_SEL_6, BUF_SEL139_6, 
        DBG_GO_2T, SPAREO2, SRAM8_WE_CLK60M_5, SRAM8_WE_CLK60M177_2, 
        BUF_SEL139_7, BUF_SEL_7, SRAM8_WE_CLK60M177_3, SPAREO3, 
        SRAM8_WE_CLK60M_4, SPAREO1_, SRAM8_WE_CLK60M_3, SPAREO4, 
        SRAM8_WE_CLK60M177_4, BUF_SEL_0, BUF_SEL2_1, BUF_SEL139_0, n312, n313, 
        n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
        n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
        n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
        n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
        n362, n363, n364, n365;
    zaoi211b SPARE_DBGFF3 ( .A(SPAREO4), .B(BUF_SEL2_0), .C(SPAREO6), .D(1'b0)
         );
    zoai21b SPARE_DBGFF4 ( .A(SPAREO0), .B(BUF_SEL_0), .C(1'b0), .Y(SPAREO9)
         );
    zoai21b SPARE_DBGFF5 ( .A(SPAREO1), .B(BUF_SEL2_1), .C(SPAREO9), .Y(
        SPAREO3) );
    zaoi211b SPARE_DBGFF2 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zdffrb SPARE_DBGFF0 ( .CK(CLK60M), .D(1'b0), .R(n323), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE_DBGFF9 ( .A(SPAREO3), .B(SPAREO6), .C(1'b0), .Y(SPAREO7) );
    zivb SPARE_DBGFF7 ( .A(SPAREO4), .Y(SPAREO5) );
    znr3b SPARE_DBGFF6 ( .A(SPAREO2), .B(BUF_SEL_1), .C(SPAREO0_), .Y(SPAREO4)
         );
    zdffrb SPARE_DBGFF1 ( .CK(CLK60M), .D(SPAREO7), .R(n323), .Q(SPAREO1), 
        .QN(SPAREO1_) );
    zivb SPARE_DBGFF8 ( .A(SPAREO5), .Y(SPAREO6) );
    zor2b U85 ( .A(BUF_SEL_4), .B(BUF_SEL_0), .Y(BUF_SEL2_0) );
    zor2b U86 ( .A(BUF_SEL_5), .B(BUF_SEL_1), .Y(BUF_SEL2_1) );
    zan2b U87 ( .A(SRAM8_WE[4]), .B(n325), .Y(SRAM8_WE_CLK60M177_4) );
    zan2b U88 ( .A(SRAM8_WE[3]), .B(n329), .Y(SRAM8_WE_CLK60M177_3) );
    zan2b U89 ( .A(SRAM8_WE[2]), .B(n328), .Y(SRAM8_WE_CLK60M177_2) );
    zan2b U90 ( .A(SRAM8_WE[7]), .B(n327), .Y(SRAM8_WE_CLK60M177_7) );
    zan2b U91 ( .A(SRAM8_WE[6]), .B(n330), .Y(SRAM8_WE_CLK60M177_6) );
    zan2b U92 ( .A(SRAM8_WE[5]), .B(n324), .Y(SRAM8_WE_CLK60M177_5) );
    zan2b U93 ( .A(SRAM8_WE[0]), .B(n331), .Y(SRAM8_WE_CLK60M177_0) );
    zan2b U94 ( .A(SRAM8_WE[1]), .B(n326), .Y(SRAM8_WE_CLK60M177_1) );
    zao21b U95 ( .A(n362), .B(n363), .C(n312), .Y(n336) );
    zivb U96 ( .A(USBPOP), .Y(n363) );
    zivb U97 ( .A(n338), .Y(n333) );
    zan2b U98 ( .A(n361), .B(BUF_SEL_7), .Y(n334) );
    zivb U99 ( .A(n336), .Y(n361) );
    znd2b U100 ( .A(n345), .B(n346), .Y(HOSTDAT[0]) );
    zaoi2x4b U101 ( .A(BUF_DAT1[24]), .B(BUF_SEL_3), .C(BUF_DAT1[16]), .D(
        BUF_SEL_2), .E(BUF_DAT1[8]), .F(BUF_SEL_1), .G(BUF_DAT1[0]), .H(n313), 
        .Y(n345) );
    zaoi2x4b U102 ( .A(BUF_DAT2[24]), .B(BUF_SEL_7), .C(BUF_DAT2[16]), .D(
        BUF_SEL_6), .E(BUF_DAT2[8]), .F(BUF_SEL_5), .G(BUF_DAT2[0]), .H(
        BUF_SEL_4), .Y(n346) );
    znd2b U103 ( .A(n347), .B(n348), .Y(HOSTDAT[1]) );
    zaoi2x4b U104 ( .A(BUF_DAT1[25]), .B(BUF_SEL_3), .C(BUF_DAT1[17]), .D(
        BUF_SEL_2), .E(BUF_DAT1[9]), .F(BUF_SEL_1), .G(BUF_DAT1[1]), .H(n313), 
        .Y(n347) );
    zaoi2x4b U105 ( .A(BUF_DAT2[25]), .B(BUF_SEL_7), .C(BUF_DAT2[17]), .D(
        BUF_SEL_6), .E(BUF_DAT2[9]), .F(BUF_SEL_5), .G(BUF_DAT2[1]), .H(
        BUF_SEL_4), .Y(n348) );
    znd2b U106 ( .A(n349), .B(n350), .Y(HOSTDAT[2]) );
    zaoi2x4b U107 ( .A(BUF_DAT1[26]), .B(BUF_SEL_3), .C(BUF_DAT1[18]), .D(
        BUF_SEL_2), .E(BUF_DAT1[10]), .F(BUF_SEL_1), .G(BUF_DAT1[2]), .H(n313), 
        .Y(n349) );
    zaoi2x4b U108 ( .A(BUF_DAT2[26]), .B(BUF_SEL_7), .C(BUF_DAT2[18]), .D(
        BUF_SEL_6), .E(BUF_DAT2[10]), .F(BUF_SEL_5), .G(BUF_DAT2[2]), .H(
        BUF_SEL_4), .Y(n350) );
    znd2b U109 ( .A(n351), .B(n352), .Y(HOSTDAT[3]) );
    zaoi2x4b U110 ( .A(BUF_DAT1[27]), .B(BUF_SEL_3), .C(BUF_DAT1[19]), .D(
        BUF_SEL_2), .E(BUF_DAT1[11]), .F(BUF_SEL_1), .G(BUF_DAT1[3]), .H(n313), 
        .Y(n351) );
    zaoi2x4b U111 ( .A(BUF_DAT2[27]), .B(BUF_SEL_7), .C(BUF_DAT2[19]), .D(
        BUF_SEL_6), .E(BUF_DAT2[11]), .F(BUF_SEL_5), .G(BUF_DAT2[3]), .H(
        BUF_SEL_4), .Y(n352) );
    znd2b U112 ( .A(n353), .B(n354), .Y(HOSTDAT[4]) );
    zaoi2x4b U113 ( .A(BUF_DAT1[28]), .B(BUF_SEL_3), .C(BUF_DAT1[20]), .D(
        BUF_SEL_2), .E(BUF_DAT1[12]), .F(BUF_SEL_1), .G(BUF_DAT1[4]), .H(n313), 
        .Y(n353) );
    zaoi2x4b U114 ( .A(BUF_DAT2[28]), .B(BUF_SEL_7), .C(BUF_DAT2[20]), .D(
        BUF_SEL_6), .E(BUF_DAT2[12]), .F(BUF_SEL_5), .G(BUF_DAT2[4]), .H(
        BUF_SEL_4), .Y(n354) );
    znd2b U115 ( .A(n355), .B(n356), .Y(HOSTDAT[5]) );
    zaoi2x4b U116 ( .A(BUF_DAT1[29]), .B(BUF_SEL_3), .C(BUF_DAT1[21]), .D(
        BUF_SEL_2), .E(BUF_DAT1[13]), .F(BUF_SEL_1), .G(BUF_DAT1[5]), .H(n313), 
        .Y(n355) );
    zaoi2x4b U117 ( .A(BUF_DAT2[29]), .B(BUF_SEL_7), .C(BUF_DAT2[21]), .D(
        BUF_SEL_6), .E(BUF_DAT2[13]), .F(BUF_SEL_5), .G(BUF_DAT2[5]), .H(
        BUF_SEL_4), .Y(n356) );
    znd2b U118 ( .A(n357), .B(n358), .Y(HOSTDAT[6]) );
    zaoi2x4b U119 ( .A(BUF_DAT1[30]), .B(BUF_SEL_3), .C(BUF_DAT1[22]), .D(
        BUF_SEL_2), .E(BUF_DAT1[14]), .F(BUF_SEL_1), .G(BUF_DAT1[6]), .H(n313), 
        .Y(n357) );
    zaoi2x4b U120 ( .A(BUF_DAT2[30]), .B(BUF_SEL_7), .C(BUF_DAT2[22]), .D(
        BUF_SEL_6), .E(BUF_DAT2[14]), .F(BUF_SEL_5), .G(BUF_DAT2[6]), .H(
        BUF_SEL_4), .Y(n358) );
    znd2b U121 ( .A(n359), .B(n360), .Y(HOSTDAT[7]) );
    zaoi2x4b U122 ( .A(BUF_SEL_3), .B(BUF_DAT1[31]), .C(BUF_SEL_2), .D(
        BUF_DAT1[23]), .E(BUF_SEL_1), .F(BUF_DAT1[15]), .G(n313), .H(BUF_DAT1
        [7]), .Y(n359) );
    zaoi2x4b U123 ( .A(BUF_SEL_7), .B(BUF_DAT2[31]), .C(BUF_SEL_6), .D(
        BUF_DAT2[23]), .E(BUF_SEL_5), .F(BUF_DAT2[15]), .G(BUF_SEL_4), .H(
        BUF_DAT2[7]), .Y(n360) );
    zao21b U124 ( .A(DI[0]), .B(n332), .C(n321), .Y(BUF_DI[0]) );
    zao21b U125 ( .A(DI[1]), .B(n332), .C(n320), .Y(BUF_DI[1]) );
    zao21b U126 ( .A(DI[2]), .B(n332), .C(n319), .Y(BUF_DI[2]) );
    zao21b U127 ( .A(DI[3]), .B(n332), .C(n318), .Y(BUF_DI[3]) );
    zao21b U128 ( .A(DI[4]), .B(n332), .C(n317), .Y(BUF_DI[4]) );
    zao21b U129 ( .A(DI[5]), .B(n332), .C(n316), .Y(BUF_DI[5]) );
    zao21b U130 ( .A(DI[6]), .B(n365), .C(n315), .Y(BUF_DI[6]) );
    zao21b U131 ( .A(DI[7]), .B(n365), .C(n314), .Y(BUF_DI[7]) );
    zao21b U132 ( .A(DI[8]), .B(n365), .C(n321), .Y(BUF_DI[8]) );
    zao21b U133 ( .A(DI[9]), .B(n365), .C(n320), .Y(BUF_DI[9]) );
    zao21b U134 ( .A(DI[10]), .B(n365), .C(n319), .Y(BUF_DI[10]) );
    zao21b U135 ( .A(DI[11]), .B(n365), .C(n318), .Y(BUF_DI[11]) );
    zao21b U136 ( .A(DI[12]), .B(n365), .C(n317), .Y(BUF_DI[12]) );
    zao21b U137 ( .A(DI[13]), .B(n365), .C(n316), .Y(BUF_DI[13]) );
    zao21b U138 ( .A(DI[14]), .B(n365), .C(n315), .Y(BUF_DI[14]) );
    zao21b U139 ( .A(DI[15]), .B(n365), .C(n314), .Y(BUF_DI[15]) );
    zao21b U140 ( .A(DI[16]), .B(n365), .C(n321), .Y(BUF_DI[16]) );
    zao21b U141 ( .A(DI[17]), .B(n365), .C(n320), .Y(BUF_DI[17]) );
    zao21b U142 ( .A(DI[18]), .B(n365), .C(n319), .Y(BUF_DI[18]) );
    zao21b U143 ( .A(DI[19]), .B(n365), .C(n318), .Y(BUF_DI[19]) );
    zao21b U144 ( .A(DI[20]), .B(n365), .C(n317), .Y(BUF_DI[20]) );
    zao21b U145 ( .A(DI[21]), .B(n365), .C(n316), .Y(BUF_DI[21]) );
    zao21b U146 ( .A(DI[22]), .B(n364), .C(n315), .Y(BUF_DI[22]) );
    zao21b U147 ( .A(DI[23]), .B(n364), .C(n314), .Y(BUF_DI[23]) );
    zao21b U148 ( .A(DI[24]), .B(n364), .C(n321), .Y(BUF_DI[24]) );
    zao21b U149 ( .A(DI[25]), .B(n364), .C(n320), .Y(BUF_DI[25]) );
    zao21b U150 ( .A(DI[26]), .B(n364), .C(n319), .Y(BUF_DI[26]) );
    zao21b U151 ( .A(DI[27]), .B(n364), .C(n318), .Y(BUF_DI[27]) );
    zao21b U152 ( .A(DI[28]), .B(n364), .C(n317), .Y(BUF_DI[28]) );
    zao21b U153 ( .A(DI[29]), .B(n364), .C(n316), .Y(BUF_DI[29]) );
    zao21b U154 ( .A(DI[30]), .B(n364), .C(n315), .Y(BUF_DI[30]) );
    zao21b U155 ( .A(DI[31]), .B(n364), .C(n314), .Y(BUF_DI[31]) );
    zao22b U156 ( .A(SRAM8_WE_CLK60M_0), .B(n332), .C(BUF_SEL_0), .D(n322), 
        .Y(BUF_WE[0]) );
    zao22b U157 ( .A(SRAM8_WE_CLK60M_1), .B(n332), .C(n322), .D(BUF_SEL_1), 
        .Y(BUF_WE[1]) );
    zao22b U158 ( .A(SRAM8_WE_CLK60M_2), .B(n332), .C(n322), .D(BUF_SEL_2), 
        .Y(BUF_WE[2]) );
    zao22b U159 ( .A(SRAM8_WE_CLK60M_3), .B(n332), .C(n322), .D(BUF_SEL_3), 
        .Y(BUF_WE[3]) );
    zao22b U160 ( .A(SRAM8_WE_CLK60M_4), .B(n332), .C(n322), .D(BUF_SEL_4), 
        .Y(BUF_WE[4]) );
    zao22b U161 ( .A(SRAM8_WE_CLK60M_5), .B(n332), .C(n322), .D(BUF_SEL_5), 
        .Y(BUF_WE[5]) );
    zao22b U162 ( .A(SRAM8_WE_CLK60M_6), .B(n332), .C(n322), .D(BUF_SEL_6), 
        .Y(BUF_WE[6]) );
    zao22b U163 ( .A(SRAM8_WE_CLK60M_7), .B(n332), .C(n322), .D(BUF_SEL_7), 
        .Y(BUF_WE[7]) );
    zivb U164 ( .A(LATCHDAT), .Y(n362) );
    zivb U165 ( .A(SRAM8_WE_CLK60M_4), .Y(n325) );
    zivb U166 ( .A(SRAM8_WE_CLK60M_3), .Y(n329) );
    zivb U167 ( .A(SRAM8_WE_CLK60M_2), .Y(n328) );
    zivb U168 ( .A(BUF_SEL_7), .Y(n344) );
    zivb U169 ( .A(BUF_SEL_6), .Y(n343) );
    zivb U170 ( .A(SRAM8_WE_CLK60M_7), .Y(n327) );
    zivb U171 ( .A(SRAM8_WE_CLK60M_6), .Y(n330) );
    zivb U172 ( .A(SRAM8_WE_CLK60M_5), .Y(n324) );
    zivb U173 ( .A(BUF_SEL_4), .Y(n341) );
    zivb U174 ( .A(BUF_SEL_5), .Y(n342) );
    zivb U175 ( .A(DBG_GO_T), .Y(n332) );
    zivb U176 ( .A(DBG_GO_T), .Y(n365) );
    zivb U177 ( .A(DBG_GO_T), .Y(n364) );
    zivb U178 ( .A(BUF_SEL_3), .Y(n340) );
    zivb U179 ( .A(SRAM8_WE_CLK60M_0), .Y(n331) );
    zivb U180 ( .A(BUF_SEL_2), .Y(n339) );
    zivb U181 ( .A(SRAM8_WE_CLK60M_1), .Y(n326) );
    zivb U182 ( .A(BUF_SEL_1), .Y(n337) );
    zivb U183 ( .A(BUF_SEL_0), .Y(n335) );
    znr2b U184 ( .A(DBG_GO_2T), .B(n332), .Y(n312) );
    znr6b U185 ( .A(BUF_SEL_6), .B(BUF_SEL_7), .C(BUF_SEL2_1), .D(BUF_SEL_2), 
        .E(BUF_SEL_3), .F(BUF_SEL_4), .Y(n313) );
    zan2b U186 ( .A(USBDAT[7]), .B(DBG_GO_T), .Y(n314) );
    zan2b U187 ( .A(USBDAT[6]), .B(DBG_GO_T), .Y(n315) );
    zan2b U188 ( .A(USBDAT[5]), .B(DBG_GO_T), .Y(n316) );
    zan2b U189 ( .A(USBDAT[4]), .B(DBG_GO_T), .Y(n317) );
    zan2b U190 ( .A(USBDAT[3]), .B(DBG_GO_T), .Y(n318) );
    zan2b U191 ( .A(USBDAT[2]), .B(DBG_GO_T), .Y(n319) );
    zan2b U192 ( .A(USBDAT[1]), .B(DBG_GO_T), .Y(n320) );
    zan2b U193 ( .A(USBDAT[0]), .B(DBG_GO_T), .Y(n321) );
    znr2b U194 ( .A(n332), .B(n362), .Y(n322) );
    zbfb U195 ( .A(HRST_), .Y(n323) );
    zdffqsb BUF_SEL_reg_0 ( .CK(CLK60M), .D(BUF_SEL139_0), .S(n323), .Q(
        BUF_SEL_0) );
    zdffqrb BUF_SEL_reg_1 ( .CK(CLK60M), .D(BUF_SEL139_1), .R(HRST_), .Q(
        BUF_SEL_1) );
    zdffqrb SRAM8_WE_CLK60M_reg_1 ( .CK(CLK60M), .D(SRAM8_WE_CLK60M177_1), .R(
        n323), .Q(SRAM8_WE_CLK60M_1) );
    zdffqrb BUF_SEL_reg_2 ( .CK(CLK60M), .D(BUF_SEL139_2), .R(HRST_), .Q(
        BUF_SEL_2) );
    zdffqrb SRAM8_WE_CLK60M_reg_0 ( .CK(CLK60M), .D(SRAM8_WE_CLK60M177_0), .R(
        HRST_), .Q(SRAM8_WE_CLK60M_0) );
    zdffqrb BUF_SEL_reg_3 ( .CK(CLK60M), .D(BUF_SEL139_3), .R(HRST_), .Q(
        BUF_SEL_3) );
    zdffqrb DBG_GO_T_reg ( .CK(CLK60M), .D(DBG_GO), .R(HRST_), .Q(DBG_GO_T) );
    zdffqrb BUF_SEL_reg_5 ( .CK(CLK60M), .D(BUF_SEL139_5), .R(HRST_), .Q(
        BUF_SEL_5) );
    zdffqrb BUF_SEL_reg_4 ( .CK(CLK60M), .D(BUF_SEL139_4), .R(HRST_), .Q(
        BUF_SEL_4) );
    zdffqrb SRAM8_WE_CLK60M_reg_5 ( .CK(CLK60M), .D(SRAM8_WE_CLK60M177_5), .R(
        HRST_), .Q(SRAM8_WE_CLK60M_5) );
    zdffqrb SRAM8_WE_CLK60M_reg_6 ( .CK(CLK60M), .D(SRAM8_WE_CLK60M177_6), .R(
        HRST_), .Q(SRAM8_WE_CLK60M_6) );
    zdffqrb SRAM8_WE_CLK60M_reg_7 ( .CK(CLK60M), .D(SRAM8_WE_CLK60M177_7), .R(
        HRST_), .Q(SRAM8_WE_CLK60M_7) );
    zdffqrb BUF_SEL_reg_6 ( .CK(CLK60M), .D(BUF_SEL139_6), .R(HRST_), .Q(
        BUF_SEL_6) );
    zdffqrb BUF_SEL_reg_7 ( .CK(CLK60M), .D(BUF_SEL139_7), .R(n323), .Q(
        BUF_SEL_7) );
    zdffqrb SRAM8_WE_CLK60M_reg_2 ( .CK(CLK60M), .D(SRAM8_WE_CLK60M177_2), .R(
        HRST_), .Q(SRAM8_WE_CLK60M_2) );
    zdffqrb DBG_GO_2T_reg ( .CK(CLK60M), .D(DBG_GO_T), .R(HRST_), .Q(DBG_GO_2T
        ) );
    zdffqrb SRAM8_WE_CLK60M_reg_3 ( .CK(CLK60M), .D(SRAM8_WE_CLK60M177_3), .R(
        HRST_), .Q(SRAM8_WE_CLK60M_3) );
    zdffqrb SRAM8_WE_CLK60M_reg_4 ( .CK(CLK60M), .D(SRAM8_WE_CLK60M177_4), .R(
        HRST_), .Q(SRAM8_WE_CLK60M_4) );
    zao211b U196 ( .A(n333), .B(BUF_SEL_0), .C(n312), .D(n334), .Y(
        BUF_SEL139_0) );
    zoai22d U197 ( .A(n335), .B(n336), .C(n337), .D(n338), .Y(BUF_SEL139_1) );
    zoai22d U198 ( .A(n337), .B(n336), .C(n339), .D(n338), .Y(BUF_SEL139_2) );
    zoai22d U199 ( .A(n339), .B(n336), .C(n340), .D(n338), .Y(BUF_SEL139_3) );
    zoai22d U200 ( .A(n340), .B(n336), .C(n341), .D(n338), .Y(BUF_SEL139_4) );
    zoai22d U201 ( .A(n341), .B(n336), .C(n342), .D(n338), .Y(BUF_SEL139_5) );
    zoai22d U202 ( .A(n342), .B(n336), .C(n343), .D(n338), .Y(BUF_SEL139_6) );
    zoai22d U203 ( .A(n343), .B(n336), .C(n344), .D(n338), .Y(BUF_SEL139_7) );
    zor3b U204 ( .A(USBPOP), .B(n312), .C(LATCHDAT), .Y(n338) );
endmodule


module DBG_BUF8X8 ( CLK, WR, DIN, DOUT1, DOUT2 );
input  [7:0] WR;
input  [31:0] DIN;
output [31:0] DOUT2;
output [31:0] DOUT1;
input  CLK;
    wire SRAM_CELL42_6__5, SRAM_CELL42_0__0, SRAM_CELL42_7__4, 
        SRAM_CELL42_1__1, SRAM_CELL42_2__4, SRAM_CELL42_4__1, SRAM_CELL42_3__5, 
        SRAM_CELL42_5__0, SRAM_CELL42_5__7, SRAM_CELL42_3__2, SRAM_CELL42_4__6, 
        SRAM_CELL42_2__3, SRAM_CELL42_1__6, SRAM_CELL42_7__3, SRAM_CELL42_0__7, 
        SRAM_CELL42_6__2, SRAM_CELL42_2__2, SRAM_CELL42_4__7, SRAM_CELL42_3__3, 
        SRAM_CELL42_5__6, SRAM_CELL42_6__3, SRAM_CELL42_0__6, SRAM_CELL42_7__2, 
        SRAM_CELL42_1__7, SRAM_CELL42_1__0, SRAM_CELL42_7__5, SRAM_CELL42_0__1, 
        SRAM_CELL42_6__4, SRAM_CELL42_5__1, SRAM_CELL42_3__4, SRAM_CELL42_4__0, 
        SRAM_CELL42_2__5, SRAM_CELL42_6__6, SRAM_CELL42_0__3, SRAM_CELL42_7__7, 
        SRAM_CELL42_1__2, SRAM_CELL42_2__7, SRAM_CELL42_4__2, SRAM_CELL42_3__6, 
        SRAM_CELL42_5__3, SRAM_CELL42_5__4, SRAM_CELL42_3__1, SRAM_CELL42_4__5, 
        SRAM_CELL42_2__0, SRAM_CELL42_1__5, SRAM_CELL42_7__0, SRAM_CELL42_0__4, 
        SRAM_CELL42_6__1, SRAM_CELL42_2__1, SRAM_CELL42_4__4, SRAM_CELL42_3__0, 
        SRAM_CELL42_5__5, SRAM_CELL42_6__0, SRAM_CELL42_0__5, SRAM_CELL42_7__1, 
        SRAM_CELL42_1__4, SRAM_CELL42_1__3, SRAM_CELL42_7__6, SRAM_CELL42_0__2, 
        SRAM_CELL42_6__7, SRAM_CELL42_5__2, SRAM_CELL42_3__7, SRAM_CELL42_4__3, 
        SRAM_CELL42_2__6;
    zmux21hb U10 ( .A(DOUT2[31]), .B(DIN[31]), .S(WR[7]), .Y(SRAM_CELL42_7__7)
         );
    zmux21hb U11 ( .A(DOUT2[30]), .B(DIN[30]), .S(WR[7]), .Y(SRAM_CELL42_7__6)
         );
    zmux21hb U12 ( .A(DOUT2[29]), .B(DIN[29]), .S(WR[7]), .Y(SRAM_CELL42_7__5)
         );
    zmux21hb U13 ( .A(DOUT2[28]), .B(DIN[28]), .S(WR[7]), .Y(SRAM_CELL42_7__4)
         );
    zmux21hb U14 ( .A(DOUT2[27]), .B(DIN[27]), .S(WR[7]), .Y(SRAM_CELL42_7__3)
         );
    zmux21hb U15 ( .A(DOUT2[26]), .B(DIN[26]), .S(WR[7]), .Y(SRAM_CELL42_7__2)
         );
    zmux21hb U16 ( .A(DOUT2[25]), .B(DIN[25]), .S(WR[7]), .Y(SRAM_CELL42_7__1)
         );
    zmux21hb U17 ( .A(DOUT2[24]), .B(DIN[24]), .S(WR[7]), .Y(SRAM_CELL42_7__0)
         );
    zmux21hb U18 ( .A(DOUT2[23]), .B(DIN[23]), .S(WR[6]), .Y(SRAM_CELL42_6__7)
         );
    zmux21hb U19 ( .A(DOUT2[22]), .B(DIN[22]), .S(WR[6]), .Y(SRAM_CELL42_6__6)
         );
    zmux21hb U20 ( .A(DOUT2[21]), .B(DIN[21]), .S(WR[6]), .Y(SRAM_CELL42_6__5)
         );
    zmux21hb U21 ( .A(DOUT2[20]), .B(DIN[20]), .S(WR[6]), .Y(SRAM_CELL42_6__4)
         );
    zmux21hb U22 ( .A(DOUT2[19]), .B(DIN[19]), .S(WR[6]), .Y(SRAM_CELL42_6__3)
         );
    zmux21hb U23 ( .A(DOUT2[18]), .B(DIN[18]), .S(WR[6]), .Y(SRAM_CELL42_6__2)
         );
    zmux21hb U24 ( .A(DOUT2[17]), .B(DIN[17]), .S(WR[6]), .Y(SRAM_CELL42_6__1)
         );
    zmux21hb U25 ( .A(DOUT2[16]), .B(DIN[16]), .S(WR[6]), .Y(SRAM_CELL42_6__0)
         );
    zmux21hb U26 ( .A(DOUT2[15]), .B(DIN[15]), .S(WR[5]), .Y(SRAM_CELL42_5__7)
         );
    zmux21hb U27 ( .A(DOUT2[14]), .B(DIN[14]), .S(WR[5]), .Y(SRAM_CELL42_5__6)
         );
    zmux21hb U28 ( .A(DOUT2[13]), .B(DIN[13]), .S(WR[5]), .Y(SRAM_CELL42_5__5)
         );
    zmux21hb U29 ( .A(DOUT2[12]), .B(DIN[12]), .S(WR[5]), .Y(SRAM_CELL42_5__4)
         );
    zmux21hb U30 ( .A(DOUT2[11]), .B(DIN[11]), .S(WR[5]), .Y(SRAM_CELL42_5__3)
         );
    zmux21hb U31 ( .A(DOUT2[10]), .B(DIN[10]), .S(WR[5]), .Y(SRAM_CELL42_5__2)
         );
    zmux21hb U32 ( .A(DOUT2[9]), .B(DIN[9]), .S(WR[5]), .Y(SRAM_CELL42_5__1)
         );
    zmux21hb U33 ( .A(DOUT2[8]), .B(DIN[8]), .S(WR[5]), .Y(SRAM_CELL42_5__0)
         );
    zmux21hb U34 ( .A(DOUT2[7]), .B(DIN[7]), .S(WR[4]), .Y(SRAM_CELL42_4__7)
         );
    zmux21hb U35 ( .A(DOUT2[6]), .B(DIN[6]), .S(WR[4]), .Y(SRAM_CELL42_4__6)
         );
    zmux21hb U36 ( .A(DOUT2[5]), .B(DIN[5]), .S(WR[4]), .Y(SRAM_CELL42_4__5)
         );
    zmux21hb U37 ( .A(DOUT2[4]), .B(DIN[4]), .S(WR[4]), .Y(SRAM_CELL42_4__4)
         );
    zmux21hb U38 ( .A(DOUT2[3]), .B(DIN[3]), .S(WR[4]), .Y(SRAM_CELL42_4__3)
         );
    zmux21hb U39 ( .A(DOUT2[2]), .B(DIN[2]), .S(WR[4]), .Y(SRAM_CELL42_4__2)
         );
    zmux21hb U40 ( .A(DOUT2[1]), .B(DIN[1]), .S(WR[4]), .Y(SRAM_CELL42_4__1)
         );
    zmux21hb U41 ( .A(DOUT2[0]), .B(DIN[0]), .S(WR[4]), .Y(SRAM_CELL42_4__0)
         );
    zmux21hb U42 ( .A(DOUT1[31]), .B(DIN[31]), .S(WR[3]), .Y(SRAM_CELL42_3__7)
         );
    zmux21hb U43 ( .A(DOUT1[30]), .B(DIN[30]), .S(WR[3]), .Y(SRAM_CELL42_3__6)
         );
    zmux21hb U44 ( .A(DOUT1[29]), .B(DIN[29]), .S(WR[3]), .Y(SRAM_CELL42_3__5)
         );
    zmux21hb U45 ( .A(DOUT1[28]), .B(DIN[28]), .S(WR[3]), .Y(SRAM_CELL42_3__4)
         );
    zmux21hb U46 ( .A(DOUT1[27]), .B(DIN[27]), .S(WR[3]), .Y(SRAM_CELL42_3__3)
         );
    zmux21hb U47 ( .A(DOUT1[26]), .B(DIN[26]), .S(WR[3]), .Y(SRAM_CELL42_3__2)
         );
    zmux21hb U48 ( .A(DOUT1[25]), .B(DIN[25]), .S(WR[3]), .Y(SRAM_CELL42_3__1)
         );
    zmux21hb U49 ( .A(DOUT1[24]), .B(DIN[24]), .S(WR[3]), .Y(SRAM_CELL42_3__0)
         );
    zmux21hb U50 ( .A(DOUT1[23]), .B(DIN[23]), .S(WR[2]), .Y(SRAM_CELL42_2__7)
         );
    zmux21hb U51 ( .A(DOUT1[22]), .B(DIN[22]), .S(WR[2]), .Y(SRAM_CELL42_2__6)
         );
    zmux21hb U52 ( .A(DOUT1[21]), .B(DIN[21]), .S(WR[2]), .Y(SRAM_CELL42_2__5)
         );
    zmux21hb U53 ( .A(DOUT1[20]), .B(DIN[20]), .S(WR[2]), .Y(SRAM_CELL42_2__4)
         );
    zmux21hb U54 ( .A(DOUT1[19]), .B(DIN[19]), .S(WR[2]), .Y(SRAM_CELL42_2__3)
         );
    zmux21hb U55 ( .A(DOUT1[18]), .B(DIN[18]), .S(WR[2]), .Y(SRAM_CELL42_2__2)
         );
    zmux21hb U56 ( .A(DOUT1[17]), .B(DIN[17]), .S(WR[2]), .Y(SRAM_CELL42_2__1)
         );
    zmux21hb U57 ( .A(DOUT1[16]), .B(DIN[16]), .S(WR[2]), .Y(SRAM_CELL42_2__0)
         );
    zmux21hb U58 ( .A(DOUT1[15]), .B(DIN[15]), .S(WR[1]), .Y(SRAM_CELL42_1__7)
         );
    zmux21hb U59 ( .A(DOUT1[14]), .B(DIN[14]), .S(WR[1]), .Y(SRAM_CELL42_1__6)
         );
    zmux21hb U60 ( .A(DOUT1[13]), .B(DIN[13]), .S(WR[1]), .Y(SRAM_CELL42_1__5)
         );
    zmux21hb U61 ( .A(DOUT1[12]), .B(DIN[12]), .S(WR[1]), .Y(SRAM_CELL42_1__4)
         );
    zmux21hb U62 ( .A(DOUT1[11]), .B(DIN[11]), .S(WR[1]), .Y(SRAM_CELL42_1__3)
         );
    zmux21hb U63 ( .A(DOUT1[10]), .B(DIN[10]), .S(WR[1]), .Y(SRAM_CELL42_1__2)
         );
    zmux21hb U64 ( .A(DOUT1[9]), .B(DIN[9]), .S(WR[1]), .Y(SRAM_CELL42_1__1)
         );
    zmux21hb U65 ( .A(DOUT1[8]), .B(DIN[8]), .S(WR[1]), .Y(SRAM_CELL42_1__0)
         );
    zmux21hb U66 ( .A(DOUT1[7]), .B(DIN[7]), .S(WR[0]), .Y(SRAM_CELL42_0__7)
         );
    zmux21hb U67 ( .A(DOUT1[6]), .B(DIN[6]), .S(WR[0]), .Y(SRAM_CELL42_0__6)
         );
    zmux21hb U68 ( .A(DOUT1[5]), .B(DIN[5]), .S(WR[0]), .Y(SRAM_CELL42_0__5)
         );
    zmux21hb U69 ( .A(DOUT1[4]), .B(DIN[4]), .S(WR[0]), .Y(SRAM_CELL42_0__4)
         );
    zmux21hb U70 ( .A(DOUT1[3]), .B(DIN[3]), .S(WR[0]), .Y(SRAM_CELL42_0__3)
         );
    zmux21hb U71 ( .A(DOUT1[2]), .B(DIN[2]), .S(WR[0]), .Y(SRAM_CELL42_0__2)
         );
    zmux21hb U72 ( .A(DOUT1[1]), .B(DIN[1]), .S(WR[0]), .Y(SRAM_CELL42_0__1)
         );
    zmux21hb U73 ( .A(DOUT1[0]), .B(DIN[0]), .S(WR[0]), .Y(SRAM_CELL42_0__0)
         );
    zdffqb SRAM_CELL_reg_7__7 ( .CK(CLK), .D(SRAM_CELL42_7__7), .Q(DOUT2[31])
         );
    zdffqb SRAM_CELL_reg_7__6 ( .CK(CLK), .D(SRAM_CELL42_7__6), .Q(DOUT2[30])
         );
    zdffqb SRAM_CELL_reg_7__5 ( .CK(CLK), .D(SRAM_CELL42_7__5), .Q(DOUT2[29])
         );
    zdffqb SRAM_CELL_reg_7__4 ( .CK(CLK), .D(SRAM_CELL42_7__4), .Q(DOUT2[28])
         );
    zdffqb SRAM_CELL_reg_7__3 ( .CK(CLK), .D(SRAM_CELL42_7__3), .Q(DOUT2[27])
         );
    zdffqb SRAM_CELL_reg_7__2 ( .CK(CLK), .D(SRAM_CELL42_7__2), .Q(DOUT2[26])
         );
    zdffqb SRAM_CELL_reg_7__1 ( .CK(CLK), .D(SRAM_CELL42_7__1), .Q(DOUT2[25])
         );
    zdffqb SRAM_CELL_reg_7__0 ( .CK(CLK), .D(SRAM_CELL42_7__0), .Q(DOUT2[24])
         );
    zdffqb SRAM_CELL_reg_6__7 ( .CK(CLK), .D(SRAM_CELL42_6__7), .Q(DOUT2[23])
         );
    zdffqb SRAM_CELL_reg_6__6 ( .CK(CLK), .D(SRAM_CELL42_6__6), .Q(DOUT2[22])
         );
    zdffqb SRAM_CELL_reg_6__5 ( .CK(CLK), .D(SRAM_CELL42_6__5), .Q(DOUT2[21])
         );
    zdffqb SRAM_CELL_reg_6__4 ( .CK(CLK), .D(SRAM_CELL42_6__4), .Q(DOUT2[20])
         );
    zdffqb SRAM_CELL_reg_6__3 ( .CK(CLK), .D(SRAM_CELL42_6__3), .Q(DOUT2[19])
         );
    zdffqb SRAM_CELL_reg_6__2 ( .CK(CLK), .D(SRAM_CELL42_6__2), .Q(DOUT2[18])
         );
    zdffqb SRAM_CELL_reg_6__1 ( .CK(CLK), .D(SRAM_CELL42_6__1), .Q(DOUT2[17])
         );
    zdffqb SRAM_CELL_reg_6__0 ( .CK(CLK), .D(SRAM_CELL42_6__0), .Q(DOUT2[16])
         );
    zdffqb SRAM_CELL_reg_5__7 ( .CK(CLK), .D(SRAM_CELL42_5__7), .Q(DOUT2[15])
         );
    zdffqb SRAM_CELL_reg_5__6 ( .CK(CLK), .D(SRAM_CELL42_5__6), .Q(DOUT2[14])
         );
    zdffqb SRAM_CELL_reg_5__5 ( .CK(CLK), .D(SRAM_CELL42_5__5), .Q(DOUT2[13])
         );
    zdffqb SRAM_CELL_reg_5__4 ( .CK(CLK), .D(SRAM_CELL42_5__4), .Q(DOUT2[12])
         );
    zdffqb SRAM_CELL_reg_5__3 ( .CK(CLK), .D(SRAM_CELL42_5__3), .Q(DOUT2[11])
         );
    zdffqb SRAM_CELL_reg_5__2 ( .CK(CLK), .D(SRAM_CELL42_5__2), .Q(DOUT2[10])
         );
    zdffqb SRAM_CELL_reg_5__1 ( .CK(CLK), .D(SRAM_CELL42_5__1), .Q(DOUT2[9])
         );
    zdffqb SRAM_CELL_reg_5__0 ( .CK(CLK), .D(SRAM_CELL42_5__0), .Q(DOUT2[8])
         );
    zdffqb SRAM_CELL_reg_4__7 ( .CK(CLK), .D(SRAM_CELL42_4__7), .Q(DOUT2[7])
         );
    zdffqb SRAM_CELL_reg_4__6 ( .CK(CLK), .D(SRAM_CELL42_4__6), .Q(DOUT2[6])
         );
    zdffqb SRAM_CELL_reg_4__5 ( .CK(CLK), .D(SRAM_CELL42_4__5), .Q(DOUT2[5])
         );
    zdffqb SRAM_CELL_reg_4__4 ( .CK(CLK), .D(SRAM_CELL42_4__4), .Q(DOUT2[4])
         );
    zdffqb SRAM_CELL_reg_4__3 ( .CK(CLK), .D(SRAM_CELL42_4__3), .Q(DOUT2[3])
         );
    zdffqb SRAM_CELL_reg_4__2 ( .CK(CLK), .D(SRAM_CELL42_4__2), .Q(DOUT2[2])
         );
    zdffqb SRAM_CELL_reg_4__1 ( .CK(CLK), .D(SRAM_CELL42_4__1), .Q(DOUT2[1])
         );
    zdffqb SRAM_CELL_reg_4__0 ( .CK(CLK), .D(SRAM_CELL42_4__0), .Q(DOUT2[0])
         );
    zdffqb SRAM_CELL_reg_3__7 ( .CK(CLK), .D(SRAM_CELL42_3__7), .Q(DOUT1[31])
         );
    zdffqb SRAM_CELL_reg_3__6 ( .CK(CLK), .D(SRAM_CELL42_3__6), .Q(DOUT1[30])
         );
    zdffqb SRAM_CELL_reg_3__5 ( .CK(CLK), .D(SRAM_CELL42_3__5), .Q(DOUT1[29])
         );
    zdffqb SRAM_CELL_reg_3__4 ( .CK(CLK), .D(SRAM_CELL42_3__4), .Q(DOUT1[28])
         );
    zdffqb SRAM_CELL_reg_3__3 ( .CK(CLK), .D(SRAM_CELL42_3__3), .Q(DOUT1[27])
         );
    zdffqb SRAM_CELL_reg_3__2 ( .CK(CLK), .D(SRAM_CELL42_3__2), .Q(DOUT1[26])
         );
    zdffqb SRAM_CELL_reg_3__1 ( .CK(CLK), .D(SRAM_CELL42_3__1), .Q(DOUT1[25])
         );
    zdffqb SRAM_CELL_reg_3__0 ( .CK(CLK), .D(SRAM_CELL42_3__0), .Q(DOUT1[24])
         );
    zdffqb SRAM_CELL_reg_2__7 ( .CK(CLK), .D(SRAM_CELL42_2__7), .Q(DOUT1[23])
         );
    zdffqb SRAM_CELL_reg_2__6 ( .CK(CLK), .D(SRAM_CELL42_2__6), .Q(DOUT1[22])
         );
    zdffqb SRAM_CELL_reg_2__5 ( .CK(CLK), .D(SRAM_CELL42_2__5), .Q(DOUT1[21])
         );
    zdffqb SRAM_CELL_reg_2__4 ( .CK(CLK), .D(SRAM_CELL42_2__4), .Q(DOUT1[20])
         );
    zdffqb SRAM_CELL_reg_2__3 ( .CK(CLK), .D(SRAM_CELL42_2__3), .Q(DOUT1[19])
         );
    zdffqb SRAM_CELL_reg_2__2 ( .CK(CLK), .D(SRAM_CELL42_2__2), .Q(DOUT1[18])
         );
    zdffqb SRAM_CELL_reg_2__1 ( .CK(CLK), .D(SRAM_CELL42_2__1), .Q(DOUT1[17])
         );
    zdffqb SRAM_CELL_reg_2__0 ( .CK(CLK), .D(SRAM_CELL42_2__0), .Q(DOUT1[16])
         );
    zdffqb SRAM_CELL_reg_1__7 ( .CK(CLK), .D(SRAM_CELL42_1__7), .Q(DOUT1[15])
         );
    zdffqb SRAM_CELL_reg_1__6 ( .CK(CLK), .D(SRAM_CELL42_1__6), .Q(DOUT1[14])
         );
    zdffqb SRAM_CELL_reg_1__5 ( .CK(CLK), .D(SRAM_CELL42_1__5), .Q(DOUT1[13])
         );
    zdffqb SRAM_CELL_reg_1__4 ( .CK(CLK), .D(SRAM_CELL42_1__4), .Q(DOUT1[12])
         );
    zdffqb SRAM_CELL_reg_1__3 ( .CK(CLK), .D(SRAM_CELL42_1__3), .Q(DOUT1[11])
         );
    zdffqb SRAM_CELL_reg_1__2 ( .CK(CLK), .D(SRAM_CELL42_1__2), .Q(DOUT1[10])
         );
    zdffqb SRAM_CELL_reg_1__1 ( .CK(CLK), .D(SRAM_CELL42_1__1), .Q(DOUT1[9])
         );
    zdffqb SRAM_CELL_reg_1__0 ( .CK(CLK), .D(SRAM_CELL42_1__0), .Q(DOUT1[8])
         );
    zdffqb SRAM_CELL_reg_0__7 ( .CK(CLK), .D(SRAM_CELL42_0__7), .Q(DOUT1[7])
         );
    zdffqb SRAM_CELL_reg_0__6 ( .CK(CLK), .D(SRAM_CELL42_0__6), .Q(DOUT1[6])
         );
    zdffqb SRAM_CELL_reg_0__5 ( .CK(CLK), .D(SRAM_CELL42_0__5), .Q(DOUT1[5])
         );
    zdffqb SRAM_CELL_reg_0__4 ( .CK(CLK), .D(SRAM_CELL42_0__4), .Q(DOUT1[4])
         );
    zdffqb SRAM_CELL_reg_0__3 ( .CK(CLK), .D(SRAM_CELL42_0__3), .Q(DOUT1[3])
         );
    zdffqb SRAM_CELL_reg_0__2 ( .CK(CLK), .D(SRAM_CELL42_0__2), .Q(DOUT1[2])
         );
    zdffqb SRAM_CELL_reg_0__1 ( .CK(CLK), .D(SRAM_CELL42_0__1), .Q(DOUT1[1])
         );
    zdffqb SRAM_CELL_reg_0__0 ( .CK(CLK), .D(SRAM_CELL42_0__0), .Q(DOUT1[0])
         );
endmodule


module UTM_DBG_MUX ( BUF_WE, UTM_WR, WE, BUF_DI, UTM_DIN, DIN, AUTOCHK, 
    BUF_OUT1, BUF_OUT2, UTM_DOUT );
input  [7:0] BUF_WE;
output [7:0] WE;
input  [31:0] BUF_OUT1;
input  [7:0] UTM_WR;
output [31:0] DIN;
input  [31:0] BUF_DI;
input  [31:0] UTM_DIN;
input  [31:0] BUF_OUT2;
output [63:0] UTM_DOUT;
input  AUTOCHK;
    wire n177, n178, n179;
    zbfb U23 ( .A(BUF_OUT1[0]), .Y(UTM_DOUT[0]) );
    zbfb U24 ( .A(BUF_OUT1[1]), .Y(UTM_DOUT[1]) );
    zbfb U25 ( .A(BUF_OUT1[2]), .Y(UTM_DOUT[2]) );
    zbfb U26 ( .A(BUF_OUT1[3]), .Y(UTM_DOUT[3]) );
    zbfb U27 ( .A(BUF_OUT1[4]), .Y(UTM_DOUT[4]) );
    zbfb U28 ( .A(BUF_OUT1[5]), .Y(UTM_DOUT[5]) );
    zbfb U29 ( .A(BUF_OUT1[6]), .Y(UTM_DOUT[6]) );
    zbfb U30 ( .A(BUF_OUT1[7]), .Y(UTM_DOUT[7]) );
    zbfb U31 ( .A(BUF_OUT1[8]), .Y(UTM_DOUT[8]) );
    zbfb U32 ( .A(BUF_OUT1[9]), .Y(UTM_DOUT[9]) );
    zbfb U33 ( .A(BUF_OUT1[10]), .Y(UTM_DOUT[10]) );
    zbfb U34 ( .A(BUF_OUT1[11]), .Y(UTM_DOUT[11]) );
    zbfb U35 ( .A(BUF_OUT1[12]), .Y(UTM_DOUT[12]) );
    zbfb U36 ( .A(BUF_OUT1[13]), .Y(UTM_DOUT[13]) );
    zbfb U37 ( .A(BUF_OUT1[14]), .Y(UTM_DOUT[14]) );
    zbfb U38 ( .A(BUF_OUT1[15]), .Y(UTM_DOUT[15]) );
    zbfb U39 ( .A(BUF_OUT1[16]), .Y(UTM_DOUT[16]) );
    zbfb U40 ( .A(BUF_OUT1[17]), .Y(UTM_DOUT[17]) );
    zbfb U41 ( .A(BUF_OUT1[18]), .Y(UTM_DOUT[18]) );
    zbfb U42 ( .A(BUF_OUT1[19]), .Y(UTM_DOUT[19]) );
    zbfb U43 ( .A(BUF_OUT1[20]), .Y(UTM_DOUT[20]) );
    zbfb U44 ( .A(BUF_OUT1[21]), .Y(UTM_DOUT[21]) );
    zbfb U45 ( .A(BUF_OUT1[22]), .Y(UTM_DOUT[22]) );
    zbfb U46 ( .A(BUF_OUT1[23]), .Y(UTM_DOUT[23]) );
    zbfb U47 ( .A(BUF_OUT1[24]), .Y(UTM_DOUT[24]) );
    zbfb U48 ( .A(BUF_OUT1[25]), .Y(UTM_DOUT[25]) );
    zbfb U49 ( .A(BUF_OUT1[26]), .Y(UTM_DOUT[26]) );
    zbfb U50 ( .A(BUF_OUT1[27]), .Y(UTM_DOUT[27]) );
    zbfb U51 ( .A(BUF_OUT1[28]), .Y(UTM_DOUT[28]) );
    zbfb U52 ( .A(BUF_OUT1[29]), .Y(UTM_DOUT[29]) );
    zbfb U53 ( .A(BUF_OUT1[30]), .Y(UTM_DOUT[30]) );
    zbfb U54 ( .A(BUF_OUT1[31]), .Y(UTM_DOUT[31]) );
    zbfb U55 ( .A(BUF_OUT2[0]), .Y(UTM_DOUT[32]) );
    zbfb U56 ( .A(BUF_OUT2[1]), .Y(UTM_DOUT[33]) );
    zbfb U57 ( .A(BUF_OUT2[2]), .Y(UTM_DOUT[34]) );
    zbfb U58 ( .A(BUF_OUT2[3]), .Y(UTM_DOUT[35]) );
    zbfb U59 ( .A(BUF_OUT2[4]), .Y(UTM_DOUT[36]) );
    zbfb U60 ( .A(BUF_OUT2[5]), .Y(UTM_DOUT[37]) );
    zbfb U61 ( .A(BUF_OUT2[6]), .Y(UTM_DOUT[38]) );
    zbfb U62 ( .A(BUF_OUT2[7]), .Y(UTM_DOUT[39]) );
    zbfb U63 ( .A(BUF_OUT2[8]), .Y(UTM_DOUT[40]) );
    zbfb U64 ( .A(BUF_OUT2[9]), .Y(UTM_DOUT[41]) );
    zbfb U65 ( .A(BUF_OUT2[10]), .Y(UTM_DOUT[42]) );
    zbfb U66 ( .A(BUF_OUT2[11]), .Y(UTM_DOUT[43]) );
    zbfb U67 ( .A(BUF_OUT2[12]), .Y(UTM_DOUT[44]) );
    zbfb U68 ( .A(BUF_OUT2[13]), .Y(UTM_DOUT[45]) );
    zbfb U69 ( .A(BUF_OUT2[14]), .Y(UTM_DOUT[46]) );
    zbfb U70 ( .A(BUF_OUT2[15]), .Y(UTM_DOUT[47]) );
    zbfb U71 ( .A(BUF_OUT2[16]), .Y(UTM_DOUT[48]) );
    zbfb U72 ( .A(BUF_OUT2[17]), .Y(UTM_DOUT[49]) );
    zbfb U73 ( .A(BUF_OUT2[18]), .Y(UTM_DOUT[50]) );
    zbfb U74 ( .A(BUF_OUT2[19]), .Y(UTM_DOUT[51]) );
    zbfb U75 ( .A(BUF_OUT2[20]), .Y(UTM_DOUT[52]) );
    zbfb U76 ( .A(BUF_OUT2[21]), .Y(UTM_DOUT[53]) );
    zbfb U77 ( .A(BUF_OUT2[22]), .Y(UTM_DOUT[54]) );
    zbfb U78 ( .A(BUF_OUT2[23]), .Y(UTM_DOUT[55]) );
    zbfb U79 ( .A(BUF_OUT2[24]), .Y(UTM_DOUT[56]) );
    zbfb U80 ( .A(BUF_OUT2[25]), .Y(UTM_DOUT[57]) );
    zbfb U81 ( .A(BUF_OUT2[26]), .Y(UTM_DOUT[58]) );
    zbfb U82 ( .A(BUF_OUT2[27]), .Y(UTM_DOUT[59]) );
    zbfb U83 ( .A(BUF_OUT2[28]), .Y(UTM_DOUT[60]) );
    zbfb U84 ( .A(BUF_OUT2[29]), .Y(UTM_DOUT[61]) );
    zbfb U85 ( .A(BUF_OUT2[30]), .Y(UTM_DOUT[62]) );
    zbfb U86 ( .A(BUF_OUT2[31]), .Y(UTM_DOUT[63]) );
    zmux21hb U87 ( .A(BUF_WE[7]), .B(UTM_WR[7]), .S(n177), .Y(WE[7]) );
    zmux21hb U88 ( .A(BUF_WE[6]), .B(UTM_WR[6]), .S(n179), .Y(WE[6]) );
    zmux21hb U89 ( .A(BUF_WE[5]), .B(UTM_WR[5]), .S(n178), .Y(WE[5]) );
    zmux21hb U90 ( .A(BUF_WE[4]), .B(UTM_WR[4]), .S(n177), .Y(WE[4]) );
    zmux21hb U91 ( .A(BUF_WE[3]), .B(UTM_WR[3]), .S(n179), .Y(WE[3]) );
    zmux21hb U92 ( .A(BUF_WE[2]), .B(UTM_WR[2]), .S(n178), .Y(WE[2]) );
    zmux21hb U93 ( .A(BUF_WE[1]), .B(UTM_WR[1]), .S(n177), .Y(WE[1]) );
    zmux21hb U94 ( .A(BUF_WE[0]), .B(UTM_WR[0]), .S(n179), .Y(WE[0]) );
    zmux21hb U95 ( .A(BUF_DI[9]), .B(UTM_DIN[9]), .S(n178), .Y(DIN[9]) );
    zmux21hb U96 ( .A(BUF_DI[8]), .B(UTM_DIN[8]), .S(n177), .Y(DIN[8]) );
    zmux21hb U97 ( .A(BUF_DI[7]), .B(UTM_DIN[7]), .S(n179), .Y(DIN[7]) );
    zmux21hb U98 ( .A(BUF_DI[6]), .B(UTM_DIN[6]), .S(n178), .Y(DIN[6]) );
    zmux21hb U99 ( .A(BUF_DI[5]), .B(UTM_DIN[5]), .S(n177), .Y(DIN[5]) );
    zmux21hb U100 ( .A(BUF_DI[4]), .B(UTM_DIN[4]), .S(n179), .Y(DIN[4]) );
    zmux21hb U101 ( .A(BUF_DI[31]), .B(UTM_DIN[31]), .S(n178), .Y(DIN[31]) );
    zmux21hb U102 ( .A(BUF_DI[30]), .B(UTM_DIN[30]), .S(n177), .Y(DIN[30]) );
    zmux21hb U103 ( .A(BUF_DI[3]), .B(UTM_DIN[3]), .S(n179), .Y(DIN[3]) );
    zmux21hb U104 ( .A(BUF_DI[29]), .B(UTM_DIN[29]), .S(n178), .Y(DIN[29]) );
    zmux21hb U105 ( .A(BUF_DI[28]), .B(UTM_DIN[28]), .S(n177), .Y(DIN[28]) );
    zmux21hb U106 ( .A(BUF_DI[27]), .B(UTM_DIN[27]), .S(n179), .Y(DIN[27]) );
    zmux21hb U107 ( .A(BUF_DI[26]), .B(UTM_DIN[26]), .S(n178), .Y(DIN[26]) );
    zmux21hb U108 ( .A(BUF_DI[25]), .B(UTM_DIN[25]), .S(n177), .Y(DIN[25]) );
    zmux21hb U109 ( .A(BUF_DI[24]), .B(UTM_DIN[24]), .S(n179), .Y(DIN[24]) );
    zmux21hb U110 ( .A(BUF_DI[23]), .B(UTM_DIN[23]), .S(n178), .Y(DIN[23]) );
    zmux21hb U111 ( .A(BUF_DI[22]), .B(UTM_DIN[22]), .S(n177), .Y(DIN[22]) );
    zmux21hb U112 ( .A(BUF_DI[21]), .B(UTM_DIN[21]), .S(n179), .Y(DIN[21]) );
    zmux21hb U113 ( .A(BUF_DI[20]), .B(UTM_DIN[20]), .S(n178), .Y(DIN[20]) );
    zmux21hb U114 ( .A(BUF_DI[2]), .B(UTM_DIN[2]), .S(n177), .Y(DIN[2]) );
    zmux21hb U115 ( .A(BUF_DI[19]), .B(UTM_DIN[19]), .S(n179), .Y(DIN[19]) );
    zmux21hb U116 ( .A(BUF_DI[18]), .B(UTM_DIN[18]), .S(n178), .Y(DIN[18]) );
    zmux21hb U117 ( .A(BUF_DI[17]), .B(UTM_DIN[17]), .S(n177), .Y(DIN[17]) );
    zmux21hb U118 ( .A(BUF_DI[16]), .B(UTM_DIN[16]), .S(n179), .Y(DIN[16]) );
    zmux21hb U119 ( .A(BUF_DI[15]), .B(UTM_DIN[15]), .S(n178), .Y(DIN[15]) );
    zmux21hb U120 ( .A(BUF_DI[14]), .B(UTM_DIN[14]), .S(n177), .Y(DIN[14]) );
    zmux21hb U121 ( .A(BUF_DI[13]), .B(UTM_DIN[13]), .S(n179), .Y(DIN[13]) );
    zmux21hb U122 ( .A(BUF_DI[12]), .B(UTM_DIN[12]), .S(n178), .Y(DIN[12]) );
    zmux21hb U123 ( .A(BUF_DI[11]), .B(UTM_DIN[11]), .S(n177), .Y(DIN[11]) );
    zmux21hb U124 ( .A(BUF_DI[10]), .B(UTM_DIN[10]), .S(n179), .Y(DIN[10]) );
    zmux21hb U125 ( .A(BUF_DI[1]), .B(UTM_DIN[1]), .S(n178), .Y(DIN[1]) );
    zmux21hb U126 ( .A(BUF_DI[0]), .B(UTM_DIN[0]), .S(n177), .Y(DIN[0]) );
    zbfh U127 ( .A(AUTOCHK), .Y(n177) );
    zbfh U128 ( .A(AUTOCHK), .Y(n178) );
    zbfh U129 ( .A(AUTOCHK), .Y(n179) );
endmodule

// USB 2.0 HS periodic FIFO control module

module HS_PER_FIFO ( ADI, USBDAT, BUISTRT, XMITSTRT, RXFIFO, LATCHDAT,
		 USBPOP, PCIWRT, PCIREAD, EOTQ, TDMAEND, RDMAEND, WPR1, WPR0,
		 UCBEO_, PCICLK, HRST_, TRST_, CLK60M, RXSTRT,
		 FFRDPCI, HOSTDAT, FCOUNT, FFULL, FEMPTY, FBE_,
		 RXPKTEND, FIFO_OK, RXERR, TEST_PACKET, TESTPKTOK,
		 SLAVEMODE, SLAVE_ACT, SLADDR, SLREAD, DATARDY, MDO,
		 BIST_RUN, BIST_RUN_C, BIST_ERR_S, ATPG_ENI,
		 BIST_PATTERN, SRAM_WR, SRAM_RUN, SRAM_ADDR, SRAM_SEL,
                 SRAM_RDATA, SRAM_ID, ATPG_CLK
	       );
input	ATPG_CLK;
input   [31:0]  BIST_PATTERN;
input   [8:0]   SRAM_ADDR;
input   [1:0]   SRAM_SEL, SRAM_ID;
input   SRAM_WR, SRAM_RUN;
output  [31:0]  SRAM_RDATA;
input	[31:0]	ADI;
input	[7:0]	USBDAT;
input	BUISTRT, XMITSTRT, RXFIFO, LATCHDAT, USBPOP, PCIWRT, PCIREAD, HRST_,
	EOTQ, TDMAEND, RDMAEND, WPR1, WPR0, PCICLK, TRST_, CLK60M, RXSTRT;
input	[3:0]	UCBEO_;
output	[31:0]	FFRDPCI;
output	[7:0]	HOSTDAT;
output	[8:0]	FCOUNT;
output	[3:0]	FBE_;
output	FFULL, FEMPTY, RXPKTEND, FIFO_OK, TESTPKTOK;
input	RXERR, TEST_PACKET, SLAVEMODE, SLAVE_ACT;
input	[7:0]	SLADDR;	// slave mode access address
input	SLREAD;		// slave mode read command queue
output	DATARDY;	// slave mode data ready
output	[31:0]	MDO;
input	BIST_RUN;	// BIST process starts
output	BIST_RUN_C;	// BIST_RUN clear
output	BIST_ERR_S;	// BIST process failed
input	ATPG_ENI;	// ATPG enable

wire [31:0] MDO, MDI, FIFO_MDI;
wire [8:0] WMA, RMA, RADDR, WADDR;
wire [3:0] TESTAD;
wire [31:0] TESTDOUT;
wire [8:0] RADDR_ATPG, WADDR_ATPG;
wire [31:0] MDI_ATPG, DOUT;

wire VDD = 1'b1;

    zbfb DNTBISTRUN ( .A(BIST_RUN), .Y(BISTRUN) );

    HS_FFCTL HS_FFCTL ( .USBDAT({USBDAT[7], USBDAT[6], USBDAT[5], USBDAT[4],
        USBDAT[3], USBDAT[2], USBDAT[1], USBDAT[0]}), .HOSTDAT({HOSTDAT[7],
        HOSTDAT[6], HOSTDAT[5], HOSTDAT[4], HOSTDAT[3], HOSTDAT[2], HOSTDAT[1]
        , HOSTDAT[0]}), .LATCHDAT(LATCHDAT), .USBPOP(USBPOP), .CLK60M(CLK60M)
        , .BUISTRT(BUISTRT), .WPR0(WPR0), .WPR1(WPR1), .EOT(EOTQ), .PCICLK(
        PCICLK), .ADI({ADI[31], ADI[30], ADI[29], ADI[28], ADI[27], ADI[26],
        ADI[25], ADI[24], ADI[23], ADI[22], ADI[21], ADI[20], ADI[19], ADI[18]
        , ADI[17], ADI[16], ADI[15], ADI[14], ADI[13], ADI[12], ADI[11],
        ADI[10], ADI[9], ADI[8], ADI[7], ADI[6], ADI[5], ADI[4], ADI[3],
        ADI[2], ADI[1], ADI[0]}), .FPUSH(FPUSH), .FPOP(FPOP), .MDO({MDO[31],
        MDO[30], MDO[29], MDO[28], MDO[27], MDO[26], MDO[25], MDO[24], MDO[23]
        , MDO[22], MDO[21], MDO[20], MDO[19], MDO[18], MDO[17], MDO[16],
        MDO[15], MDO[14], MDO[13], MDO[12], MDO[11], MDO[10], MDO[9], MDO[8],
        MDO[7], MDO[6], MDO[5], MDO[4], MDO[3], MDO[2], MDO[1], MDO[0]}),
        .MDI(FIFO_MDI), .WMA(WMA),
        .RMA({RMA[8], RMA[7], RMA[6], RMA[5], RMA[4]
        , RMA[3], RMA[2], RMA[1], RMA[0]}), .PCIWRT(PCIWRT), .PCIREAD(PCIREAD)
        , .RXFIFO(RXFIFO), .UCBEO_({UCBEO_[3], UCBEO_[2], UCBEO_[1], UCBEO_[0]
        }), .RXSTRT(RXSTRT), .XMITSTRT(XMITSTRT), .FIFO_OK(FIFO_OK), .FFRDPCI(
        {FFRDPCI[31], FFRDPCI[30], FFRDPCI[29], FFRDPCI[28], FFRDPCI[27],
        FFRDPCI[26], FFRDPCI[25], FFRDPCI[24], FFRDPCI[23], FFRDPCI[22],
        FFRDPCI[21], FFRDPCI[20], FFRDPCI[19], FFRDPCI[18], FFRDPCI[17],
        FFRDPCI[16], FFRDPCI[15], FFRDPCI[14], FFRDPCI[13], FFRDPCI[12],
        FFRDPCI[11], FFRDPCI[10], FFRDPCI[9], FFRDPCI[8], FFRDPCI[7],
        FFRDPCI[6], FFRDPCI[5], FFRDPCI[4], FFRDPCI[3], FFRDPCI[2], FFRDPCI[1]
        , FFRDPCI[0]}), .FBE_({FBE_[3], FBE_[2], FBE_[1], FBE_[0]}), .RDMAEND(
        //RDMAEND), .RXPKTEND(RXPKTEND), .HRST_(HRST_), .FCOUNT({FCOUNT[8],
        RDMAEND), .RXPKTEND(RXPKTEND), .TRST_(TRST_), .FCOUNT({FCOUNT[8],
        FCOUNT[7], FCOUNT[6], FCOUNT[5], FCOUNT[4], FCOUNT[3], FCOUNT[2],
        FCOUNT[1], FCOUNT[0]}), .FFULL(FFULL), .FEMPTY(FEMPTY),
	.TDMAEND(TDMAEND), .RXERR(RXERR), .TEST_PACKET(TEST_PACKET),
	.TESTAD(TESTAD), .TESTDOUT(TESTDOUT), .TESTPKTOK(TESTPKTOK),
	.ATPG_ENI(ATPG_ENI) );

    TESTDATA TESTDATA ( .PCICLK(PCICLK), .TEST_PACKET(TEST_PACKET),
        .TESTAD(TESTAD), .TESTDOUT(TESTDOUT) );

    HS_ACCESS HS_ACCESS ( .SLADDR(SLADDR), .SLREAD(SLREAD), .RMA(RMA),
	.RADDR(RADDR), .SLAVEMODE(SLAVEMODE), .DATARDY(DATARDY),
	.FPOP(FPOP), .RD(RD), .PCICLK(PCICLK), .TRST_(TRST_),
	.SLAVE_ACT(SLAVE_ACT), .FPUSH(FPUSH), .WR(WR), .MDO(MDO),
	.BIST_RUN(BISTRUN), .BIST_RUN_C(BIST_RUN_C), .FIFO_MDI(FIFO_MDI),
	.MDI(MDI), .WMA(WMA), .WADDR(WADDR), .BIST_ERR_S(BIST_ERR_S),
	.RADDR_ATPG(RADDR_ATPG), .WADDR_ATPG(WADDR_ATPG),
	.MDI_ATPG(MDI_ATPG), .ASYNCFIFO(1'b0),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_ID(SRAM_ID), .SRAM_WR(SRAM_WR),
        .SRAM_RUN(SRAM_RUN), .SRAM_RDATA(SRAM_RDATA),
	.ATPG_CLK(ATPG_CLK) );

    FIFO_ATPG_MUX FIFO_ATPG_MUX ( .ATPG_ENI(ATPG_ENI), .DOUT(DOUT),
	.MDI_ATPG(MDI_ATPG), .MDO(MDO) );

    //ssram260x32 ssram260x32 ( .RCLK(PCICLK), .WCLK(PCICLK),
    dpram260x32 dpram260x32 ( .RCLK(PCICLK), .WCLK(PCICLK),
	.WR(WR), .RD(RD), .DIN31(MDI[31]), .DIN30(MDI[30]),
	.DIN29(MDI[29]), .DIN28(MDI[28]), .DIN27(MDI[27]), .DIN26(MDI[26]),
	.DIN25(MDI[25]), .DIN24(MDI[24]), .DIN23(MDI[23]), .DIN22(MDI[22]),
	.DIN21(MDI[21]), .DIN20(MDI[20]), .DIN19(MDI[19]), .DIN18(MDI[18]),
	.DIN17(MDI[17]), .DIN16(MDI[16]), .DIN15(MDI[15]), .DIN14(MDI[14]),
	.DIN13(MDI[13]), .DIN12(MDI[12]), .DIN11(MDI[11]), .DIN10(MDI[10]),
	.DIN9(MDI[9]), .DIN8(MDI[8]), .DIN7(MDI[7]), .DIN6(MDI[6]),
	.DIN5(MDI[5]), .DIN4(MDI[4]), .DIN3(MDI[3]), .DIN2(MDI[2]),
	.DIN1(MDI[1]), .DIN0(MDI[0]),
	.DOUT31(DOUT[31]), .DOUT30(DOUT[30]), .DOUT29(DOUT[29]),
	.DOUT28(DOUT[28]), .DOUT27(DOUT[27]), .DOUT26(DOUT[26]),
        .DOUT25(DOUT[25]), .DOUT24(DOUT[24]), .DOUT23(DOUT[23]),
	.DOUT22(DOUT[22]), .DOUT21(DOUT[21]), .DOUT20(DOUT[20]),
	.DOUT19(DOUT[19]), .DOUT18(DOUT[18]), .DOUT17(DOUT[17]),
	.DOUT16(DOUT[16]), .DOUT15(DOUT[15]), .DOUT14(DOUT[14]),
        .DOUT13(DOUT[13]), .DOUT12(DOUT[12]), .DOUT11(DOUT[11]),
	.DOUT10(DOUT[10]), .DOUT9(DOUT[9]), .DOUT8(DOUT[8]),
	.DOUT7(DOUT[7]), .DOUT6(DOUT[6]), .DOUT5(DOUT[5]),
	.DOUT4(DOUT[4]), .DOUT3(DOUT[3]), .DOUT2(DOUT[2]),
        .DOUT1(DOUT[1]), .DOUT0(DOUT[0]),
	.RADDR8(RADDR[8]), .RADDR7(RADDR[7]), .RADDR6(RADDR[6]),
	.RADDR5(RADDR[5]), .RADDR4(RADDR[4]), .RADDR3(RADDR[3]),
	.RADDR2(RADDR[2]), .RADDR1(RADDR[1]), .RADDR0(RADDR[0]),
	.WADDR8(WADDR[8]), .WADDR7(WADDR[7]), .WADDR6(WADDR[6]),
	.WADDR5(WADDR[5]), .WADDR4(WADDR[4]), .WADDR3(WADDR[3]),
	.WADDR2(WADDR[2]), .WADDR1(WADDR[1]), .WADDR0(WADDR[0]),
	.RESET(HRST_) );


    /*ssram260x32 ssram260x32 ( .DOUT(MDO), .DIN(MDI), .WADDR(WADDR),
        .RADDR(RADDR), .WR(WR), .RD(RD), .RCLK(PCICLK), .WCLK(PCICLK),
	.RESET(HRST_) );*/

    /*ssram512x32 ssram512x32 ( .DOUT(MDO), .DIN(MDI), .WADDR(WMA),
        .RADDR(RMA), .WR(FPUSH), .RD(FPOP), .RCLK(PCICLK), .WCLK(PCICLK),
	.RESET(VDD) );*/

    /*ssram512x32 ssram512x32 ( .MDO31(MDO[31]), .MDO30(MDO[30]), .MDO29(MDO[29]
        ), .MDO28(MDO[28]), .MDO27(MDO[27]), .MDO26(MDO[26]), .MDO25(MDO[25])
        , .MDO24(MDO[24]), .MDO23(MDO[23]), .MDO22(MDO[22]), .MDO21(MDO[21]),
        .MDO20(MDO[20]), .MDO19(MDO[19]), .MDO18(MDO[18]), .MDO17(MDO[17]),
        .MDO16(MDO[16]), .MDO15(MDO[15]), .MDO14(MDO[14]), .MDO13(MDO[13]),
        .MDO12(MDO[12]), .MDO11(MDO[11]), .MDO10(MDO[10]), .MDO9(MDO[9]),
        .MDO8(MDO[8]), .MDO7(MDO[7]), .MDO6(MDO[6]), .MDO5(MDO[5]), .MDO4(
        MDO[4]), .MDO3(MDO[3]), .MDO2(MDO[2]), .MDO1(MDO[1]), .MDO0(MDO[0]),
        .MDI31(MDI[31]), .MDI30(MDI[30]), .MDI29(MDI[29]), .MDI28(MDI[28]),
        .MDI27(MDI[27]), .MDI26(MDI[26]), .MDI25(MDI[25]), .MDI24(MDI[24]),
        .MDI23(MDI[23]), .MDI22(MDI[22]), .MDI21(MDI[21]), .MDI20(MDI[20]),
        .MDI19(MDI[19]), .MDI18(MDI[18]), .MDI17(MDI[17]), .MDI16(MDI[16]),
        .MDI15(MDI[15]), .MDI14(MDI[14]), .MDI13(MDI[13]), .MDI12(MDI[12]),
        .MDI11(MDI[11]), .MDI10(MDI[10]), .MDI9(MDI[9]), .MDI8(MDI[8]), .MDI7(
        MDI[7]), .MDI6(MDI[6]), .MDI5(MDI[5]), .MDI4(MDI[4]), .MDI3(MDI[3]),
        .MDI2(MDI[2]), .MDI1(MDI[1]), .MDI0(MDI[0]), .WMA8(WMA[8]), .WMA7(
        WMA[7]), .WMA6(WMA[6]), .WMA5(WMA[5]), .WMA4(WMA[4]), .WMA3(WMA[3]),
        .WMA2(WMA[2]), .WMA1(WMA[1]), .WMA0(WMA[0]), .RMA8(RMA[8]), .RMA7(
        RMA[7]), .RMA6(RMA[6]), .RMA5(RMA[5]), .RMA4(RMA[4]), .RMA3(RMA[3]),
        .RMA2(RMA[2]), .RMA1(RMA[1]), .RMA0(RMA[0]), .WR(FPUSH), .RD(FPOP),
        .CLK(PCICLK), .RAMRSTZ(VDD) );*/

endmodule

// USB 2.0 HS asynchronous FIFO control module

module HS_ASYNC_FIFO ( ADI, USBDAT, BUISTRT, XMITSTRT, RXFIFO, LATCHDAT,
		 USBPOP, PCIWRT, PCIREAD, EOTQ, TDMAEND, RDMAEND, WPR1, WPR0,
		 UCBEO_, PCICLK, HRST_, TRST_, CLK60M, RXSTRT,
		 FFRDPCI, HOSTDAT, FCOUNT, FFULL, FEMPTY, FBE_,
		 RXPKTEND, FIFO_OK, RXERR, TEST_PACKET, TESTPKTOK,
		 SLAVEMODE, SLAVE_ACT, SLADDR, SLREAD, DATARDY, MDO,
		 BIST_RUN, BIST_RUN_C, BIST_ERR_S, ATPG_ENI,
		 BIST_PATTERN, SRAM_WR, SRAM_RUN, SRAM_ADDR, SRAM_SEL,
                 SRAM_RDATA, SRAM_ID, ATPG_CLK
	       );
input	ATPG_CLK;
input   [31:0]  BIST_PATTERN;
input   [8:0]   SRAM_ADDR;
input   [1:0]   SRAM_SEL, SRAM_ID;
input   SRAM_WR, SRAM_RUN;
output  [31:0]  SRAM_RDATA;
input	[31:0]	ADI;
input	[7:0]	USBDAT;
input	BUISTRT, XMITSTRT, RXFIFO, LATCHDAT, USBPOP, PCIWRT, PCIREAD, HRST_,
	EOTQ, TDMAEND, RDMAEND, WPR1, WPR0, PCICLK, TRST_, CLK60M, RXSTRT;
input	[3:0]	UCBEO_;
output	[31:0]	FFRDPCI;
output	[7:0]	HOSTDAT;
output	[8:0]	FCOUNT;
output	[3:0]	FBE_;
output	FFULL, FEMPTY, RXPKTEND, FIFO_OK, TESTPKTOK;
input	RXERR, TEST_PACKET, SLAVEMODE, SLAVE_ACT;
input	[7:0]	SLADDR;	// slave mode access address
input	SLREAD;		// slave mode read command queue
output	DATARDY;	// slave mode data ready
output	[31:0]	MDO;
input	BIST_RUN;	// BIST process starts
output	BIST_RUN_C;	// BIST_RUN clear
output	BIST_ERR_S;	// BIST process failed
input	ATPG_ENI;	// ATPG enable

wire [31:0] MDO, MDI, FIFO_MDI;
wire [8:0] WMA, RMA, RADDR, WADDR;
wire [3:0] TESTAD;
wire [31:0] TESTDOUT;
wire [8:0] RADDR_ATPG, WADDR_ATPG;
wire [31:0] MDI_ATPG, DOUT;

wire VDD = 1'b1;

    zbfb DNTBISTRUN ( .A(BIST_RUN), .Y(BISTRUN) );

    HS_FFCTL HS_FFCTL ( .USBDAT({USBDAT[7], USBDAT[6], USBDAT[5], USBDAT[4],
        USBDAT[3], USBDAT[2], USBDAT[1], USBDAT[0]}), .HOSTDAT({HOSTDAT[7],
        HOSTDAT[6], HOSTDAT[5], HOSTDAT[4], HOSTDAT[3], HOSTDAT[2], HOSTDAT[1]
        , HOSTDAT[0]}), .LATCHDAT(LATCHDAT), .USBPOP(USBPOP), .CLK60M(CLK60M)
        , .BUISTRT(BUISTRT), .WPR0(WPR0), .WPR1(WPR1), .EOT(EOTQ), .PCICLK(
        PCICLK), .ADI({ADI[31], ADI[30], ADI[29], ADI[28], ADI[27], ADI[26],
        ADI[25], ADI[24], ADI[23], ADI[22], ADI[21], ADI[20], ADI[19], ADI[18]
        , ADI[17], ADI[16], ADI[15], ADI[14], ADI[13], ADI[12], ADI[11],
        ADI[10], ADI[9], ADI[8], ADI[7], ADI[6], ADI[5], ADI[4], ADI[3],
        ADI[2], ADI[1], ADI[0]}), .FPUSH(FPUSH), .FPOP(FPOP), .MDO({MDO[31],
        MDO[30], MDO[29], MDO[28], MDO[27], MDO[26], MDO[25], MDO[24], MDO[23]
        , MDO[22], MDO[21], MDO[20], MDO[19], MDO[18], MDO[17], MDO[16],
        MDO[15], MDO[14], MDO[13], MDO[12], MDO[11], MDO[10], MDO[9], MDO[8],
        MDO[7], MDO[6], MDO[5], MDO[4], MDO[3], MDO[2], MDO[1], MDO[0]}),
        .MDI(FIFO_MDI), .WMA(WMA),
        .RMA({RMA[8], RMA[7], RMA[6], RMA[5], RMA[4]
        , RMA[3], RMA[2], RMA[1], RMA[0]}), .PCIWRT(PCIWRT), .PCIREAD(PCIREAD)
        , .RXFIFO(RXFIFO), .UCBEO_({UCBEO_[3], UCBEO_[2], UCBEO_[1], UCBEO_[0]
        }), .RXSTRT(RXSTRT), .XMITSTRT(XMITSTRT), .FIFO_OK(FIFO_OK), .FFRDPCI(
        {FFRDPCI[31], FFRDPCI[30], FFRDPCI[29], FFRDPCI[28], FFRDPCI[27],
        FFRDPCI[26], FFRDPCI[25], FFRDPCI[24], FFRDPCI[23], FFRDPCI[22],
        FFRDPCI[21], FFRDPCI[20], FFRDPCI[19], FFRDPCI[18], FFRDPCI[17],
        FFRDPCI[16], FFRDPCI[15], FFRDPCI[14], FFRDPCI[13], FFRDPCI[12],
        FFRDPCI[11], FFRDPCI[10], FFRDPCI[9], FFRDPCI[8], FFRDPCI[7],
        FFRDPCI[6], FFRDPCI[5], FFRDPCI[4], FFRDPCI[3], FFRDPCI[2], FFRDPCI[1]
        , FFRDPCI[0]}), .FBE_({FBE_[3], FBE_[2], FBE_[1], FBE_[0]}), .RDMAEND(
        //RDMAEND), .RXPKTEND(RXPKTEND), .HRST_(HRST_), .FCOUNT({FCOUNT[8],
        RDMAEND), .RXPKTEND(RXPKTEND), .TRST_(TRST_), .FCOUNT({FCOUNT[8],
        FCOUNT[7], FCOUNT[6], FCOUNT[5], FCOUNT[4], FCOUNT[3], FCOUNT[2],
        FCOUNT[1], FCOUNT[0]}), .FFULL(FFULL), .FEMPTY(FEMPTY),
	.TDMAEND(TDMAEND), .RXERR(RXERR), .TEST_PACKET(TEST_PACKET),
	.TESTAD(TESTAD), .TESTDOUT(TESTDOUT), .TESTPKTOK(TESTPKTOK),
	.ATPG_ENI(ATPG_ENI) );

    TESTDATA TESTDATA ( .PCICLK(PCICLK), .TEST_PACKET(TEST_PACKET),
        .TESTAD(TESTAD), .TESTDOUT(TESTDOUT) );

    HS_ACCESS HS_ACCESS ( .SLADDR(SLADDR), .SLREAD(SLREAD), .RMA(RMA),
	.RADDR(RADDR), .SLAVEMODE(SLAVEMODE), .DATARDY(DATARDY),
	.FPOP(FPOP), .RD(RD), .PCICLK(PCICLK), .TRST_(TRST_),
	.SLAVE_ACT(SLAVE_ACT), .FPUSH(FPUSH), .WR(WR), .MDO(MDO),
	.BIST_RUN(BISTRUN), .BIST_RUN_C(BIST_RUN_C), .FIFO_MDI(FIFO_MDI),
	.MDI(MDI), .WMA(WMA), .WADDR(WADDR), .BIST_ERR_S(BIST_ERR_S),
	.RADDR_ATPG(RADDR_ATPG), .WADDR_ATPG(WADDR_ATPG),
	.MDI_ATPG(MDI_ATPG), .ASYNCFIFO(1'b1),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_ID(SRAM_ID), .SRAM_WR(SRAM_WR),
        .SRAM_RUN(SRAM_RUN), .SRAM_RDATA(SRAM_RDATA),
	.ATPG_CLK(ATPG_CLK) );

    FIFO_ATPG_MUX FIFO_ATPG_MUX ( .ATPG_ENI(ATPG_ENI), .DOUT(DOUT),
	.MDI_ATPG(MDI_ATPG), .MDO(MDO) );

    //ssram132x32 ssram132x32 ( .RCLK(PCICLK), .WCLK(PCICLK),
    dpram132x32 dpram132x32 ( .RCLK(PCICLK), .WCLK(PCICLK),
	.WR(WR), .RD(RD), .DIN31(MDI[31]), .DIN30(MDI[30]),
	.DIN29(MDI[29]), .DIN28(MDI[28]), .DIN27(MDI[27]), .DIN26(MDI[26]),
	.DIN25(MDI[25]), .DIN24(MDI[24]), .DIN23(MDI[23]), .DIN22(MDI[22]),
	.DIN21(MDI[21]), .DIN20(MDI[20]), .DIN19(MDI[19]), .DIN18(MDI[18]),
	.DIN17(MDI[17]), .DIN16(MDI[16]), .DIN15(MDI[15]), .DIN14(MDI[14]),
	.DIN13(MDI[13]), .DIN12(MDI[12]), .DIN11(MDI[11]), .DIN10(MDI[10]),
	.DIN9(MDI[9]), .DIN8(MDI[8]), .DIN7(MDI[7]), .DIN6(MDI[6]),
	.DIN5(MDI[5]), .DIN4(MDI[4]), .DIN3(MDI[3]), .DIN2(MDI[2]),
	.DIN1(MDI[1]), .DIN0(MDI[0]),
	.DOUT31(DOUT[31]), .DOUT30(DOUT[30]), .DOUT29(DOUT[29]),
	.DOUT28(DOUT[28]), .DOUT27(DOUT[27]), .DOUT26(DOUT[26]),
        .DOUT25(DOUT[25]), .DOUT24(DOUT[24]), .DOUT23(DOUT[23]),
	.DOUT22(DOUT[22]), .DOUT21(DOUT[21]), .DOUT20(DOUT[20]),
	.DOUT19(DOUT[19]), .DOUT18(DOUT[18]), .DOUT17(DOUT[17]),
	.DOUT16(DOUT[16]), .DOUT15(DOUT[15]), .DOUT14(DOUT[14]),
        .DOUT13(DOUT[13]), .DOUT12(DOUT[12]), .DOUT11(DOUT[11]),
	.DOUT10(DOUT[10]), .DOUT9(DOUT[9]), .DOUT8(DOUT[8]),
	.DOUT7(DOUT[7]), .DOUT6(DOUT[6]), .DOUT5(DOUT[5]),
	.DOUT4(DOUT[4]), .DOUT3(DOUT[3]), .DOUT2(DOUT[2]),
        .DOUT1(DOUT[1]), .DOUT0(DOUT[0]),
	/*.RADDR8(RADDR[8]),*/ .RADDR7(RADDR[7]), .RADDR6(RADDR[6]),
	.RADDR5(RADDR[5]), .RADDR4(RADDR[4]), .RADDR3(RADDR[3]),
	.RADDR2(RADDR[2]), .RADDR1(RADDR[1]), .RADDR0(RADDR[0]),
	/*.WADDR8(WADDR[8]),*/ .WADDR7(WADDR[7]), .WADDR6(WADDR[6]),
	.WADDR5(WADDR[5]), .WADDR4(WADDR[4]), .WADDR3(WADDR[3]),
	.WADDR2(WADDR[2]), .WADDR1(WADDR[1]), .WADDR0(WADDR[0]),
	.RESET(HRST_) );

endmodule

// USB 2.0 HS DEBUG_PORT FIFO control module

module DBG_FIFO (   DBG_BUF_WE, DI,
                    DBGPORT_BUF1, DBGPORT_BUF2,
                    DBG_GO,
                    LATCHDAT, USBPOP, USBDAT, HOSTDAT,
		    UTM_WR, UTM_DIN, UTM_DOUT, AUTOCHK,
                    CLK60M, HRST_ );
input	[7:0]	UTM_WR;
input	[31:0]	UTM_DIN;
output	[63:0]	UTM_DOUT;
input	AUTOCHK;
input   [7:0]   DBG_BUF_WE;
input   [31:0]  DI;
output  [31:0]  DBGPORT_BUF1, DBGPORT_BUF2;
input   DBG_GO;
input   LATCHDAT, USBPOP;
input   [7:0]   USBDAT;
output  [7:0]   HOSTDAT;
input   CLK60M, HRST_;

wire  [31:0]  BUF_DI, DIN;
wire  [7:0]   BUF_WE, WE;

    DBG_FFCTL DBG_FFCTL ( .SRAM8_WE(DBG_BUF_WE), .DI(DI),
	.BUF_WE(BUF_WE), .BUF_DI(BUF_DI), .BUF_DAT1(DBGPORT_BUF1),
	.BUF_DAT2(DBGPORT_BUF2), .DBG_GO(DBG_GO),
	.LATCHDAT(LATCHDAT), .USBPOP(USBPOP), .USBDAT(USBDAT),
	.HOSTDAT(HOSTDAT), .CLK60M(CLK60M), .HRST_(HRST_) );

    UTM_DBG_MUX UTM_DBG_MUX ( .BUF_WE(BUF_WE), .UTM_WR(UTM_WR),
	.WE(WE), .BUF_DI(BUF_DI), .UTM_DIN(UTM_DIN), .DIN(DIN),
	.BUF_OUT1(DBGPORT_BUF1), .BUF_OUT2(DBGPORT_BUF2),
	.UTM_DOUT(UTM_DOUT), .AUTOCHK(AUTOCHK) );

    DBG_BUF8X8 DBG_BUF8X8 ( .CLK(CLK60M), .WR(WE), .DIN(DIN),
	.DOUT1(DBGPORT_BUF1), .DOUT2(DBGPORT_BUF2) );

endmodule


module HS_BMUSM ( HCIGNT, FIFOGNT, RDMAEND, TDMAEND, TXREQ, RXREQ, RFREQ_S, 
    RFLUSH_S, EOTQ, XMITSTRT, TXTHRESH, XMITNULL, BUFEND, MABORTS, TABORTR, 
    BUSTMOUT, FEMPTY, MYPMACK, RXSTRT, QRXERR, RXTHRESH, RXPKTEND, BUSFREE, 
    UGNTI_, HCIREQ, PCICLK, HRST_, DISTXDLY, EOF, DISTXDLY2, BMUSM_RST_EN, 
    DBUFERR, DISPFIFO, ZEROLEN, DISRXZERO, BUI_GO, DISPFIFO2, ENBMUSMRST, 
    DMA_IDLE, ATPG_ENI, FIFO_OK );
input  EOTQ, XMITSTRT, TXTHRESH, XMITNULL, BUFEND, MABORTS, TABORTR, BUSTMOUT, 
    FEMPTY, MYPMACK, RXSTRT, QRXERR, RXTHRESH, RXPKTEND, BUSFREE, UGNTI_, 
    HCIREQ, PCICLK, HRST_, DISTXDLY, EOF, DISTXDLY2, BMUSM_RST_EN, DBUFERR, 
    DISPFIFO, ZEROLEN, DISRXZERO, BUI_GO, DISPFIFO2, ENBMUSMRST, ATPG_ENI, 
    FIFO_OK;
output HCIGNT, FIFOGNT, RDMAEND, TDMAEND, TXREQ, RXREQ, RFREQ_S, RFLUSH_S, 
    DMA_IDLE;
    wire TXFFPR_2, SPAREO6, TXFFNX_2, ownc0, SPAREO0_, SPAREO8, SPAREO1, 
        RXFFNX_2, SPAREO9, FIFOREQ, RXFFPR_2, SPAREO0, SPAREO7, ownc1, 
        TXFFPR_1, SPAREO5, TXFFNX_1, ownd1, TXRST_, RXFFNX_0, SPAREO2, 
        RXFFPR_0, RXFFNX_1, ownd0, SPAREO3, SPAREO1_, RXFFPR_1, TXFFPR_0, 
        SPAREO4, TXFFNX_0, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
        n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
        n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
        n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
        n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
        n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
        n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233;
    zoai21b SPARE715 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE712 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zaoi211b SPARE713 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zoai21b SPARE714 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    znr3b SPARE716 ( .A(SPAREO2), .B(FIFOREQ), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE718 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE711 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    znd3b SPARE719 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE710 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE717 ( .A(SPAREO4), .Y(SPAREO5) );
    zivb U324 ( .A(DISPFIFO2), .Y(n1214) );
    zivb U325 ( .A(DISTXDLY), .Y(n1194) );
    zan2b U326 ( .A(TXTHRESH), .B(n1197), .Y(n1218) );
    zivb U327 ( .A(FEMPTY), .Y(n1201) );
    zan3b U328 ( .A(n1204), .B(n1205), .C(n1206), .Y(n1203) );
    zivb U329 ( .A(ZEROLEN), .Y(n1228) );
    zor2b U330 ( .A(FEMPTY), .B(n1200), .Y(n1233) );
    zivb U331 ( .A(RXTHRESH), .Y(n1206) );
    zor2b U332 ( .A(RXPKTEND), .B(n1211), .Y(n1204) );
    znd2b U333 ( .A(BUSTMOUT), .B(MYPMACK), .Y(n1212) );
    zan3b U334 ( .A(n1189), .B(n1190), .C(BUSFREE), .Y(n1188) );
    zor2b U335 ( .A(RXFFPR_2), .B(n1224), .Y(n1225) );
    zivb U336 ( .A(n1225), .Y(n1205) );
    zivb U337 ( .A(TXTHRESH), .Y(n1182) );
    zan3b U338 ( .A(BUFEND), .B(n1232), .C(TXFFPR_1), .Y(n1183) );
    zor2b U339 ( .A(TABORTR), .B(MABORTS), .Y(n1179) );
    zivb U340 ( .A(n1211), .Y(n1175) );
    zivb U341 ( .A(DISPFIFO), .Y(n1222) );
    zao32b U342 ( .A(TXREQ), .B(n1198), .C(n1202), .D(TDMAEND), .E(TXFFPR_0), 
        .Y(n1176) );
    zivb U343 ( .A(BUFEND), .Y(n1198) );
    zan2b U344 ( .A(n1232), .B(n1219), .Y(n1177) );
    zan2b U345 ( .A(n1200), .B(RXFFPR_1), .Y(n1207) );
    zmux31hb U346 ( .A(RXFFPR_1), .B(RXFFPR_0), .D0(n1229), .D1(RXTHRESH), 
        .D2(n1179), .Y(n1208) );
    zivb U347 ( .A(n1204), .Y(n1200) );
    zivb U348 ( .A(n1179), .Y(n1202) );
    zmux21lb U349 ( .A(n1230), .B(n1231), .S(RXFFPR_0), .Y(n1187) );
    zan3b U350 ( .A(n1189), .B(n1192), .C(BUSFREE), .Y(n1172) );
    zivb U351 ( .A(UGNTI_), .Y(n1189) );
    zivb U352 ( .A(HCIREQ), .Y(n1221) );
    zor2b U353 ( .A(TXREQ), .B(RXREQ), .Y(FIFOREQ) );
    zivb U354 ( .A(FIFOREQ), .Y(n1191) );
    znr5b U355 ( .A(RXFFPR_0), .B(n1169), .C(RXFFPR_2), .D(TXFFPR_1), .E(
        RXFFPR_1), .Y(DMA_IDLE) );
    zor2b U356 ( .A(TXFFPR_0), .B(TXFFPR_2), .Y(n1169) );
    zivb U357 ( .A(n1169), .Y(n1232) );
    zivb U358 ( .A(n1227), .Y(RFLUSH_S) );
    zivb U359 ( .A(n1226), .Y(RFREQ_S) );
    zor2b U360 ( .A(n1220), .B(n1225), .Y(n1226) );
    zivb U361 ( .A(n1223), .Y(RDMAEND) );
    zor2b U362 ( .A(RXFFPR_1), .B(n1209), .Y(n1223) );
    zdffqrb TXFFPR_reg_2 ( .CK(PCICLK), .D(TXFFNX_2), .R(TXRST_), .Q(TXFFPR_2)
         );
    zivb U363 ( .A(TXFFPR_2), .Y(n1178) );
    zdffqrb TXFFPR_reg_1 ( .CK(PCICLK), .D(TXFFNX_1), .R(TXRST_), .Q(TXFFPR_1)
         );
    zivb U364 ( .A(TXFFPR_1), .Y(n1219) );
    zdffrb TXFFPR_reg_0 ( .CK(PCICLK), .D(TXFFNX_0), .R(TXRST_), .Q(TXFFPR_0), 
        .QN(n1197) );
    zdffqrb RXFFPR_reg_2 ( .CK(PCICLK), .D(RXFFNX_2), .R(TXRST_), .Q(RXFFPR_2)
         );
    zivb U365 ( .A(RXFFPR_2), .Y(n1209) );
    zdffqrb RXFFPR_reg_1 ( .CK(PCICLK), .D(RXFFNX_1), .R(TXRST_), .Q(RXFFPR_1)
         );
    zivb U366 ( .A(RXFFPR_1), .Y(n1224) );
    zdffqrb RXFFPR_reg_0 ( .CK(PCICLK), .D(RXFFNX_0), .R(TXRST_), .Q(RXFFPR_0)
         );
    zivb U367 ( .A(RXFFPR_0), .Y(n1220) );
    zdffrb ownc0_reg ( .CK(PCICLK), .D(ownd0), .R(HRST_), .Q(ownc0), .QN(n1190
        ) );
    zdffrb ownc1_reg ( .CK(PCICLK), .D(ownd1), .R(HRST_), .Q(ownc1), .QN(n1192
        ) );
    zan3b U368 ( .A(RXFFPR_0), .B(n1209), .C(FIFO_OK), .Y(RXREQ) );
    znr3b U369 ( .A(TXFFPR_2), .B(n1197), .C(n1219), .Y(TXREQ) );
    znr2b U370 ( .A(ownc0), .B(n1192), .Y(HCIGNT) );
    znr2b U371 ( .A(ownc1), .B(n1190), .Y(FIFOGNT) );
    znr2b U372 ( .A(TXFFPR_1), .B(n1178), .Y(TDMAEND) );
    znr3b U373 ( .A(n1220), .B(n1223), .C(n1211), .Y(n1167) );
    zmux21hb U374 ( .A(n1217), .B(n1218), .S(TXFFPR_1), .Y(n1168) );
    zao211b U375 ( .A(DISPFIFO2), .B(n1170), .C(ATPG_ENI), .D(n1171), .Y(
        TXRST_) );
    zoa21d U376 ( .A(n1172), .B(n1173), .C(FIFOREQ), .Y(ownd0) );
    zoa21d U377 ( .A(n1174), .B(HCIGNT), .C(HCIREQ), .Y(ownd1) );
    zao222b U378 ( .A(n1175), .B(n1176), .C(n1177), .D(XMITSTRT), .E(n1168), 
        .F(n1178), .Y(TXFFNX_0) );
    zao21b U379 ( .A(TXREQ), .B(n1179), .C(n1180), .Y(TXFFNX_1) );
    zao222b U380 ( .A(n1175), .B(n1181), .C(TXREQ), .D(n1179), .E(n1182), .F(
        n1183), .Y(TXFFNX_2) );
    zor3b U381 ( .A(n1167), .B(n1184), .C(n1185), .Y(RXFFNX_2) );
    zor3b U382 ( .A(n1167), .B(n1186), .C(n1187), .Y(RXFFNX_0) );
    zoa21d U383 ( .A(n1188), .B(FIFOGNT), .C(n1191), .Y(n1174) );
    zoa21d U384 ( .A(BMUSM_RST_EN), .B(DISTXDLY2), .C(n1194), .Y(n1193) );
    znr2d U385 ( .A(BUI_GO), .B(n1195), .Y(n1171) );
    zoa211b U386 ( .A(n1175), .B(n1197), .C(TXFFPR_1), .D(n1198), .Y(n1196) );
    zoa21d U387 ( .A(n1196), .B(n1168), .C(n1178), .Y(n1180) );
    zoa21d U388 ( .A(n1200), .B(n1201), .C(n1202), .Y(n1199) );
    zoa21d U389 ( .A(n1203), .B(RFLUSH_S), .C(FEMPTY), .Y(n1184) );
    zoa21d U390 ( .A(n1207), .B(n1208), .C(n1209), .Y(RXFFNX_1) );
    zoa22b U391 ( .A(RXFFPR_2), .B(n1200), .C(RXFFPR_1), .D(n1211), .Y(n1210)
         );
    zan4b U392 ( .A(n1200), .B(RFREQ_S), .C(n1202), .D(n1212), .Y(n1186) );
    zan2d U393 ( .A(HRST_), .B(n1214), .Y(n1213) );
    zmux21hd U394 ( .A(n1216), .B(EOF), .S(n1193), .Y(n1215) );
    zivf U395 ( .A(HRST_), .Y(n1216) );
    zao21b U396 ( .A(DBUFERR), .B(n1222), .C(EOTQ), .Y(n1211) );
    zor3b U397 ( .A(RXFFPR_2), .B(RXFFPR_1), .C(n1220), .Y(n1227) );
    zmux21ld U398 ( .A(n1213), .B(n1170), .S(ENBMUSMRST), .Y(n1195) );
    zinr2b U399 ( .A(TXFFPR_0), .B(XMITNULL), .Y(n1217) );
    zoa21d U400 ( .A(DISRXZERO), .B(n1228), .C(RXSTRT), .Y(n1229) );
    zao21b U401 ( .A(HCIGNT), .B(n1221), .C(FIFOGNT), .Y(n1173) );
    zoai22b U402 ( .A(n1202), .B(n1227), .C(n1199), .D(n1226), .Y(n1185) );
    zao21b U403 ( .A(TXREQ), .B(BUFEND), .C(TDMAEND), .Y(n1181) );
    zivf U404 ( .A(n1215), .Y(n1170) );
    zor3b U405 ( .A(n1179), .B(n1210), .C(FEMPTY), .Y(n1231) );
    zao21b U406 ( .A(n1233), .B(n1206), .C(n1225), .Y(n1230) );
endmodule


module HS_BMUTM ( WPR, TFCOMPL, RFCOMPL, BUSTMOUT, BUFEND, BCNT10, BCNT9, 
    BCNT8, BCNT7, BCNT6, BCNT5, BCNT4, BCNT3, BCNT2, BCNT1, BCNT0, TFGNT, 
    RFGNT, BCNTBT40, UMORE, UMORE2LN, MBE3_, MBE2_, MBE1_, MBE0_, BUFPTR1, 
    BUFPTR2, MAXLEN, RFREQ_S, TXREQ, RFLUSH_S, FEMPTY, FIFOGNT, PMSTR, RDYACK, 
    NEARFEMP, WPRLD, TXFIFO, RXFIFO, FCFG, FBE_, PCICLK, HRST_, BOUNDRY, 
    BOUNDRY_T, DIS_BURST, HCIGNT );
output [31:0] WPR;
input  [31:0] BUFPTR2;
input  [3:0] FBE_;
input  [31:0] BUFPTR1;
input  [10:0] MAXLEN;
input  RFREQ_S, TXREQ, RFLUSH_S, FEMPTY, FIFOGNT, PMSTR, RDYACK, NEARFEMP, 
    WPRLD, TXFIFO, RXFIFO, FCFG, PCICLK, HRST_, DIS_BURST, HCIGNT;
output TFCOMPL, RFCOMPL, BUSTMOUT, BUFEND, BCNT10, BCNT9, BCNT8, BCNT7, BCNT6, 
    BCNT5, BCNT4, BCNT3, BCNT2, BCNT1, BCNT0, TFGNT, RFGNT, BCNTBT40, UMORE, 
    UMORE2LN, MBE3_, MBE2_, MBE1_, MBE0_, BOUNDRY, BOUNDRY_T;
    wire BUFPTR2_LT_17, WPR387_4, BUFPTR2_LT_7, WPR387_17, SPAREO6, WPR387_30, 
        WPR_NX_21, BCNT_NX_2, BCNT462_5, BUFPTR2_LT363_17, BTIMER304_1, 
        BUFPTR2_LT363_2, BTIMER290_1, BTIMER_1, WPR_NX_14, WPR387_22, 
        WPR_NX_28, WPR_NX_6, BUFPTR2_LT363_19, WPR387_25, NEARBEND, WPR_NX_1, 
        SPAREO0_, BUFPTR2_LT_9, BOUNDRY_T425, WPR387_19, WPR_NX_13, SPAREO8, 
        BCNT_NX_5, BUFPTR2_LT_19, BUFPTR2_LT363_5, BUFPTR2_LT363_10, BCNT462_2, 
        BCNT_NX_10, WPR_NX_26, WPR_NX_8, SPAREO1, WPR387_10, BUFPTR2_LT_0, 
        BUFPTR2_LT_10, WPR387_3, BUFPTR2_LT_18, BUFPTR2_LT363_4, BUFPTR2_LT_8, 
        WPR_NX_12, SPAREO9, WPR387_18, BCNT_NX_4, WPR387_24, WPR_NX_0, 
        BUFPTR2_LT363_18, BUFPTR2_LT_11, WPR387_2, WPR387_11, BUFPTR2_LT_1, 
        SPAREO0, WPR_NX_27, WPR_NX_9, BUFPTR2_LT363_11, BCNT462_3, BCNT462_4, 
        BUFPTR2_LT363_16, WPR_NX_20, BUFPTR2_LT_6, SPAREO7, WPR387_16, 
        WPR387_31, BUFPTR2_LT_16, WPR387_5, SIZEB4, WPR_NX_29, WPR387_23, 
        WPR_NX_7, BCNT_NX_3, BTIMER_0, WPR_NX_15, BTIMER304_0, BUFPTR2_LT363_3, 
        WPR387_7, BUFPTR2_LT363_8, BUFPTR2_LT_14, BCNT_NX_8, BUFPTR2_LT_4, 
        WPR387_14, SPAREO5, WPR_NX_22, WPR387_28, BUFPTR2_LT363_14, BCNT462_6, 
        BTIMER304_2, BUFPTR2_LT363_1, WPR_NX_17, BTIMER_2, BCNT_NX_1, 
        WPR_NX_30, BTIMER290_2, WPR_NX_5, WPR387_21, BCNT462_10, BCNT462_8, 
        WPR_NX_2, BCNTBT20, BCNT_NX_6, WPR387_26, WPR_NX_10, WPR387_9, 
        BUFPTR2_LT363_6, BUFPTR2_LT363_13, BCNT462_1, WPR_NX_25, BTIMER_4, 
        WPR_NX_19, SPAREO2, WPR387_13, BUFPTR2_LT_3, WPR387_0, BUFPTR2_LT_13, 
        WPR387_8, BTIMER304_4, BUFPTR2_LT363_7, BCNT_NX_7, WPR_NX_11, 
        BTIMER290_4, WPR_NX_3, WPR387_27, BCNT462_9, WPR387_1, BUFPTR2_LT_12, 
        WPR387_12, WPR_NX_18, SPAREO3, BUFPTR2_LT_2, SPAREO1_, WPR_NX_24, 
        BCNT462_0, BUFPTR2_LT363_12, BUFPTR2_LT363_15, BCNT462_7, WPR387_29, 
        WPR_NX_23, BCNT_NX_9, BUFPTR2_LT_5, SPAREO4, WPR387_15, WPR387_6, 
        BUFPTR2_LT363_9, BUFPTR2_LT_15, WPR_NX_4, WPR387_20, WPR_NX_16, 
        BTIMER_3, BCNT_NX_0, WPR_NX_31, BTIMER290_3, BTIMER304_3, 
        BUFPTR2_LT363_0, n593, n594, n595, n596, n597, n598, n599, n600, n601, 
        n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, 
        n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, 
        n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, 
        n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, 
        n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, 
        n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, 
        n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, 
        n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, 
        n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, 
        n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, 
        n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, 
        n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
        n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, 
        n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, 
        n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, 
        n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, 
        n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, 
        n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, 
        n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
        n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, 
        n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, 
        n854;
    zoai21b SPARE715 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zaoi211b SPARE712 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zaoi211b SPARE713 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zoai21b SPARE714 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    znr3b SPARE716 ( .A(SPAREO2), .B(TFCOMPL), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE718 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE711 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    znd3b SPARE719 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE710 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    zivb SPARE717 ( .A(SPAREO4), .Y(SPAREO5) );
    znd2b U202 ( .A(WPR[25]), .B(WPR[23]), .Y(n653) );
    znd2b U203 ( .A(WPR[22]), .B(WPR[24]), .Y(n651) );
    znd2b U204 ( .A(WPR[9]), .B(WPR[8]), .Y(n655) );
    znd2b U205 ( .A(WPR[7]), .B(WPR[6]), .Y(n656) );
    znd3b U206 ( .A(WPR[3]), .B(WPR[4]), .C(WPR[5]), .Y(n657) );
    zan2b U207 ( .A(n597), .B(n786), .Y(n780) );
    zan3b U208 ( .A(MBE0_), .B(MBE2_), .C(n792), .Y(n791) );
    znd2b U209 ( .A(n779), .B(n810), .Y(n732) );
    znr2b U210 ( .A(BCNT5), .B(BCNT4), .Y(n737) );
    znd2b U211 ( .A(WPR[29]), .B(WPR[30]), .Y(n650) );
    znd3b U212 ( .A(WPR[27]), .B(WPR[28]), .C(WPR[26]), .Y(n679) );
    znd2b U213 ( .A(WPR[27]), .B(WPR[26]), .Y(n722) );
    znr2b U214 ( .A(n651), .B(n653), .Y(n652) );
    znd3b U215 ( .A(WPR[24]), .B(WPR[23]), .C(WPR[22]), .Y(n713) );
    znd2b U216 ( .A(WPR[22]), .B(WPR[23]), .Y(n725) );
    znd2b U217 ( .A(WPR[19]), .B(WPR[20]), .Y(n684) );
    znd2b U218 ( .A(WPR[21]), .B(WPR[18]), .Y(n683) );
    zan2b U219 ( .A(WPR[18]), .B(WPR[19]), .Y(n675) );
    zan2b U220 ( .A(WPR[14]), .B(WPR[15]), .Y(n672) );
    zor2b U221 ( .A(n693), .B(n692), .Y(n694) );
    znd2b U222 ( .A(WPR[12]), .B(WPR[11]), .Y(n693) );
    znd2b U223 ( .A(WPR[10]), .B(WPR[13]), .Y(n692) );
    zivb U224 ( .A(n694), .Y(n673) );
    zan2b U225 ( .A(WPR[10]), .B(WPR[11]), .Y(n670) );
    zor2b U226 ( .A(n615), .B(n644), .Y(n614) );
    zivb U227 ( .A(n690), .Y(n615) );
    znr3b U228 ( .A(n657), .B(n656), .C(n655), .Y(n690) );
    zan2b U229 ( .A(WPR[7]), .B(WPR[6]), .Y(n698) );
    znr2b U230 ( .A(n658), .B(n701), .Y(n699) );
    znd2b U231 ( .A(WPR[3]), .B(WPR[4]), .Y(n658) );
    znd2b U232 ( .A(WPR[2]), .B(n784), .Y(n644) );
    zivd U233 ( .A(n784), .Y(n740) );
    znd2b U234 ( .A(WPR[1]), .B(n779), .Y(n648) );
    zivd U235 ( .A(n779), .Y(n741) );
    ziv11b U236 ( .A(RDYACK), .Y(n620), .Z(n619) );
    znd2b U237 ( .A(n784), .B(n627), .Y(n728) );
    zivb U238 ( .A(n738), .Y(n749) );
    znr3b U239 ( .A(BCNT9), .B(BCNT7), .C(BCNT3), .Y(n765) );
    znr2b U240 ( .A(BCNT4), .B(BCNT8), .Y(n766) );
    znr2b U241 ( .A(BCNT5), .B(BCNT10), .Y(n767) );
    znr2b U242 ( .A(BCNT6), .B(BCNT2), .Y(n768) );
    znd2b U243 ( .A(BTIMER_3), .B(n601), .Y(n638) );
    znd2b U244 ( .A(n728), .B(n733), .Y(n746) );
    zivb U245 ( .A(n729), .Y(n745) );
    znd2b U246 ( .A(n732), .B(n731), .Y(n744) );
    zivc U247 ( .A(n750), .Y(n736) );
    znd2b U248 ( .A(BCNT0), .B(n742), .Y(n759) );
    zivb U249 ( .A(n782), .Y(n742) );
    znd2b U250 ( .A(n758), .B(n757), .Y(BCNT_NX_8) );
    znd2b U251 ( .A(BCNT8), .B(n754), .Y(n757) );
    znd2b U252 ( .A(n754), .B(n753), .Y(BCNT_NX_7) );
    znd2b U253 ( .A(BCNT7), .B(n756), .Y(n753) );
    znd2b U254 ( .A(BCNT6), .B(n763), .Y(n755) );
    znd2b U255 ( .A(BTIMER_1), .B(BTIMER_0), .Y(n641) );
    zivb U256 ( .A(n679), .Y(n642) );
    znd2b U257 ( .A(n617), .B(WPR[26]), .Y(n666) );
    znr2b U258 ( .A(n726), .B(n725), .Y(n727) );
    zivf U259 ( .A(n682), .Y(n676) );
    zivb U260 ( .A(n674), .Y(n671) );
    znd2b U261 ( .A(n671), .B(WPR[14]), .Y(n662) );
    znd2b U262 ( .A(n605), .B(WPR[12]), .Y(n661) );
    znd2b U263 ( .A(n700), .B(n699), .Y(n716) );
    zivc U264 ( .A(n716), .Y(n697) );
    znd2b U265 ( .A(n603), .B(WPR[4]), .Y(n668) );
    zivb U266 ( .A(n700), .Y(n706) );
    znd2b U267 ( .A(n645), .B(n644), .Y(n705) );
    zivb U268 ( .A(n646), .Y(n704) );
    znd2b U269 ( .A(n649), .B(n648), .Y(n660) );
    znd2b U270 ( .A(WPR[0]), .B(n782), .Y(n720) );
    znr2b U271 ( .A(n782), .B(WPR[0]), .Y(n719) );
    znd2b U272 ( .A(n762), .B(n761), .Y(BCNT_NX_4) );
    znd2b U273 ( .A(n736), .B(n734), .Y(n762) );
    znd2b U274 ( .A(BCNT4), .B(n750), .Y(n761) );
    zivb U275 ( .A(n762), .Y(n764) );
    zivb U276 ( .A(n733), .Y(n748) );
    zan3b U277 ( .A(WPR[9]), .B(WPR[11]), .C(WPR[3]), .Y(n820) );
    zor2b U278 ( .A(n805), .B(n811), .Y(n823) );
    zor2b U279 ( .A(WPR[0]), .B(n817), .Y(n826) );
    zmux21lb U280 ( .A(n812), .B(n811), .S(n593), .Y(n821) );
    zor2b U281 ( .A(n813), .B(n814), .Y(n812) );
    zivb U282 ( .A(n817), .Y(n813) );
    znr2b U283 ( .A(BCNT7), .B(BCNT9), .Y(n635) );
    znr2b U284 ( .A(BCNT5), .B(BCNT10), .Y(n637) );
    znd3b U285 ( .A(n623), .B(n622), .C(n621), .Y(n629) );
    znr2b U286 ( .A(n628), .B(n627), .Y(n630) );
    znr2b U287 ( .A(BCNT1), .B(BCNT0), .Y(n628) );
    znd3b U288 ( .A(n626), .B(n624), .C(n625), .Y(n631) );
    znr2b U289 ( .A(BCNT7), .B(BCNT3), .Y(n626) );
    znr2b U290 ( .A(BCNT4), .B(BCNT8), .Y(n625) );
    zivb U291 ( .A(n819), .Y(n789) );
    znr5b U292 ( .A(n620), .B(MBE3_), .C(HCIGNT), .D(n769), .E(n770), .Y(
        BOUNDRY_T425) );
    zivb U293 ( .A(PMSTR), .Y(n769) );
    zivb U294 ( .A(n770), .Y(BOUNDRY) );
    znd8b U295 ( .A(WPR[5]), .B(WPR[8]), .C(WPR[7]), .D(WPR[4]), .E(WPR[6]), 
        .F(WPR[2]), .G(WPR[10]), .H(n820), .Y(n770) );
    zao22b U296 ( .A(FBE_[0]), .B(n596), .C(TFGNT), .D(n775), .Y(MBE0_) );
    zivb U297 ( .A(MBE0_), .Y(n785) );
    zan2b U298 ( .A(n814), .B(n811), .Y(n774) );
    zivb U299 ( .A(n815), .Y(n814) );
    zivb U300 ( .A(MBE1_), .Y(n786) );
    zmux21lb U301 ( .A(n822), .B(n823), .S(WPR[1]), .Y(n773) );
    zao22b U302 ( .A(FBE_[3]), .B(n596), .C(TFGNT), .D(n772), .Y(MBE3_) );
    zivb U303 ( .A(MBE3_), .Y(n818) );
    zan2b U304 ( .A(BCNTBT40), .B(TFGNT), .Y(UMORE2LN) );
    zan2b U305 ( .A(BCNTBT20), .B(TFGNT), .Y(UMORE) );
    znd3b U306 ( .A(n633), .B(n634), .C(n632), .Y(BCNTBT40) );
    znr2b U307 ( .A(BCNT7), .B(BCNT9), .Y(n633) );
    znr2b U308 ( .A(BCNT10), .B(BCNT6), .Y(n632) );
    zivb U309 ( .A(n816), .Y(RFGNT) );
    zor2b U310 ( .A(n804), .B(n808), .Y(n816) );
    zivb U311 ( .A(RXFIFO), .Y(n808) );
    zivb U312 ( .A(n805), .Y(TFGNT) );
    zor2b U313 ( .A(n803), .B(n804), .Y(n805) );
    zivb U314 ( .A(TXFIFO), .Y(n803) );
    zivb U315 ( .A(FIFOGNT), .Y(n804) );
    znr6b U316 ( .A(n776), .B(BCNT1), .C(BCNT0), .D(BCNT3), .E(BCNT4), .F(
        BCNT2), .Y(BUFEND) );
    zan3b U317 ( .A(n599), .B(n639), .C(n771), .Y(BUSTMOUT) );
    zan2b U318 ( .A(RXFIFO), .B(n778), .Y(RFCOMPL) );
    zao32b U319 ( .A(RFLUSH_S), .B(n825), .C(NEARFEMP), .D(RFREQ_S), .E(n777), 
        .Y(n778) );
    zivb U320 ( .A(FEMPTY), .Y(n825) );
    znr3b U321 ( .A(n631), .B(n630), .C(n629), .Y(NEARBEND) );
    zivb U322 ( .A(BCNT8), .Y(n735) );
    zdffqrb BTIMER_reg_3 ( .CK(PCICLK), .D(BTIMER304_3), .R(HRST_), .Q(
        BTIMER_3) );
    zdffqrb BTIMER_reg_1 ( .CK(PCICLK), .D(BTIMER304_1), .R(HRST_), .Q(
        BTIMER_1) );
    zivb U323 ( .A(BTIMER_1), .Y(n806) );
    zdffb BUFPTR2_LT_reg_19 ( .CK(PCICLK), .D(BUFPTR2_LT363_19), .Q(
        BUFPTR2_LT_19), .QN(n801) );
    zdffqb BUFPTR2_LT_reg_18 ( .CK(PCICLK), .D(BUFPTR2_LT363_18), .Q(
        BUFPTR2_LT_18) );
    zdffqb BUFPTR2_LT_reg_17 ( .CK(PCICLK), .D(BUFPTR2_LT363_17), .Q(
        BUFPTR2_LT_17) );
    zdffqb BUFPTR2_LT_reg_16 ( .CK(PCICLK), .D(BUFPTR2_LT363_16), .Q(
        BUFPTR2_LT_16) );
    zdffqb BUFPTR2_LT_reg_15 ( .CK(PCICLK), .D(BUFPTR2_LT363_15), .Q(
        BUFPTR2_LT_15) );
    zdffqb BUFPTR2_LT_reg_14 ( .CK(PCICLK), .D(BUFPTR2_LT363_14), .Q(
        BUFPTR2_LT_14) );
    zdffqb BUFPTR2_LT_reg_13 ( .CK(PCICLK), .D(BUFPTR2_LT363_13), .Q(
        BUFPTR2_LT_13) );
    zdffqb BUFPTR2_LT_reg_12 ( .CK(PCICLK), .D(BUFPTR2_LT363_12), .Q(
        BUFPTR2_LT_12) );
    zdffqb BUFPTR2_LT_reg_11 ( .CK(PCICLK), .D(BUFPTR2_LT363_11), .Q(
        BUFPTR2_LT_11) );
    zdffqb BUFPTR2_LT_reg_10 ( .CK(PCICLK), .D(BUFPTR2_LT363_10), .Q(
        BUFPTR2_LT_10) );
    zdffqb BUFPTR2_LT_reg_9 ( .CK(PCICLK), .D(BUFPTR2_LT363_9), .Q(
        BUFPTR2_LT_9) );
    zdffqb BUFPTR2_LT_reg_8 ( .CK(PCICLK), .D(BUFPTR2_LT363_8), .Q(
        BUFPTR2_LT_8) );
    zdffqb BUFPTR2_LT_reg_7 ( .CK(PCICLK), .D(BUFPTR2_LT363_7), .Q(
        BUFPTR2_LT_7) );
    zdffqb BUFPTR2_LT_reg_6 ( .CK(PCICLK), .D(BUFPTR2_LT363_6), .Q(
        BUFPTR2_LT_6) );
    zdffqb BUFPTR2_LT_reg_5 ( .CK(PCICLK), .D(BUFPTR2_LT363_5), .Q(
        BUFPTR2_LT_5) );
    zdffqb BUFPTR2_LT_reg_4 ( .CK(PCICLK), .D(BUFPTR2_LT363_4), .Q(
        BUFPTR2_LT_4) );
    zdffqb BUFPTR2_LT_reg_3 ( .CK(PCICLK), .D(BUFPTR2_LT363_3), .Q(
        BUFPTR2_LT_3) );
    zdffqb BUFPTR2_LT_reg_2 ( .CK(PCICLK), .D(BUFPTR2_LT363_2), .Q(
        BUFPTR2_LT_2) );
    zdffqb BUFPTR2_LT_reg_1 ( .CK(PCICLK), .D(BUFPTR2_LT363_1), .Q(
        BUFPTR2_LT_1) );
    zdffqb BUFPTR2_LT_reg_0 ( .CK(PCICLK), .D(BUFPTR2_LT363_0), .Q(
        BUFPTR2_LT_0) );
    zdffqrb WPR_reg_31 ( .CK(PCICLK), .D(WPR387_31), .R(HRST_), .Q(WPR[31]) );
    zdffqrb WPR_reg_30 ( .CK(PCICLK), .D(WPR387_30), .R(HRST_), .Q(WPR[30]) );
    zdffqrb WPR_reg_29 ( .CK(PCICLK), .D(WPR387_29), .R(HRST_), .Q(WPR[29]) );
    zivb U324 ( .A(WPR[29]), .Y(n678) );
    zdffqrb WPR_reg_28 ( .CK(PCICLK), .D(WPR387_28), .R(HRST_), .Q(WPR[28]) );
    zdffqrb WPR_reg_27 ( .CK(PCICLK), .D(WPR387_27), .R(HRST_), .Q(WPR[27]) );
    zivb U325 ( .A(WPR[27]), .Y(n680) );
    zdffqrb WPR_reg_26 ( .CK(PCICLK), .D(WPR387_26), .R(HRST_), .Q(WPR[26]) );
    zdffqrb WPR_reg_25 ( .CK(PCICLK), .D(WPR387_25), .R(HRST_), .Q(WPR[25]) );
    zdffqrb WPR_reg_24 ( .CK(PCICLK), .D(WPR387_24), .R(HRST_), .Q(WPR[24]) );
    zdffqrb WPR_reg_23 ( .CK(PCICLK), .D(WPR387_23), .R(HRST_), .Q(WPR[23]) );
    zdffqrb WPR_reg_22 ( .CK(PCICLK), .D(WPR387_22), .R(HRST_), .Q(WPR[22]) );
    zivb U326 ( .A(WPR[22]), .Y(n711) );
    zdffqrb WPR_reg_21 ( .CK(PCICLK), .D(WPR387_21), .R(HRST_), .Q(WPR[21]) );
    zivb U327 ( .A(WPR[21]), .Y(n685) );
    zdffqrb WPR_reg_20 ( .CK(PCICLK), .D(WPR387_20), .R(HRST_), .Q(WPR[20]) );
    zdffqrb WPR_reg_19 ( .CK(PCICLK), .D(WPR387_19), .R(HRST_), .Q(WPR[19]) );
    zivb U328 ( .A(WPR[19]), .Y(n687) );
    zdffqrb WPR_reg_18 ( .CK(PCICLK), .D(WPR387_18), .R(HRST_), .Q(WPR[18]) );
    zivb U329 ( .A(WPR[18]), .Y(n686) );
    zdffqrb WPR_reg_17 ( .CK(PCICLK), .D(WPR387_17), .R(HRST_), .Q(WPR[17]) );
    zivb U330 ( .A(WPR[17]), .Y(n688) );
    zdffqrb WPR_reg_16 ( .CK(PCICLK), .D(WPR387_16), .R(HRST_), .Q(WPR[16]) );
    zdffqrb WPR_reg_15 ( .CK(PCICLK), .D(WPR387_15), .R(HRST_), .Q(WPR[15]) );
    zivb U331 ( .A(WPR[15]), .Y(n691) );
    zdffqrb WPR_reg_14 ( .CK(PCICLK), .D(WPR387_14), .R(HRST_), .Q(WPR[14]) );
    zivb U332 ( .A(WPR[14]), .Y(n689) );
    zdffqrb WPR_reg_13 ( .CK(PCICLK), .D(WPR387_13), .R(HRST_), .Q(WPR[13]) );
    zivb U333 ( .A(WPR[13]), .Y(n695) );
    zdffqrb WPR_reg_12 ( .CK(PCICLK), .D(WPR387_12), .R(HRST_), .Q(WPR[12]) );
    zdffqrb WPR_reg_11 ( .CK(PCICLK), .D(WPR387_11), .R(HRST_), .Q(WPR[11]) );
    zdffqrb WPR_reg_10 ( .CK(PCICLK), .D(WPR387_10), .R(HRST_), .Q(WPR[10]) );
    zivb U334 ( .A(WPR[10]), .Y(n709) );
    zdffqrb WPR_reg_9 ( .CK(PCICLK), .D(WPR387_9), .R(HRST_), .Q(WPR[9]) );
    zivb U335 ( .A(WPR[9]), .Y(n696) );
    zdffqrb WPR_reg_8 ( .CK(PCICLK), .D(WPR387_8), .R(HRST_), .Q(WPR[8]) );
    zdffqrb WPR_reg_7 ( .CK(PCICLK), .D(WPR387_7), .R(HRST_), .Q(WPR[7]) );
    zdffqrb WPR_reg_6 ( .CK(PCICLK), .D(WPR387_6), .R(HRST_), .Q(WPR[6]) );
    zivb U336 ( .A(WPR[6]), .Y(n717) );
    zdffqrb WPR_reg_5 ( .CK(PCICLK), .D(WPR387_5), .R(HRST_), .Q(WPR[5]) );
    zivb U337 ( .A(WPR[5]), .Y(n701) );
    zdffqrb WPR_reg_4 ( .CK(PCICLK), .D(WPR387_4), .R(HRST_), .Q(WPR[4]) );
    zdffqrb WPR_reg_3 ( .CK(PCICLK), .D(WPR387_3), .R(HRST_), .Q(WPR[3]) );
    zivb U338 ( .A(WPR[3]), .Y(n707) );
    zdffqrb WPR_reg_2 ( .CK(PCICLK), .D(WPR387_2), .R(HRST_), .Q(WPR[2]) );
    zivb U339 ( .A(WPR[2]), .Y(n702) );
    zdffqrb WPR_reg_1 ( .CK(PCICLK), .D(WPR387_1), .R(HRST_), .Q(WPR[1]) );
    zivb U340 ( .A(WPR[1]), .Y(n703) );
    zdffqrb WPR_reg_0 ( .CK(PCICLK), .D(WPR387_0), .R(HRST_), .Q(WPR[0]) );
    zivb U341 ( .A(WPR[0]), .Y(n811) );
    zdffrb BCNT_reg_10 ( .CK(PCICLK), .D(BCNT462_10), .R(HRST_), .Q(BCNT10), 
        .QN(n623) );
    zdffqrb BCNT_reg_4 ( .CK(PCICLK), .D(BCNT462_4), .R(HRST_), .Q(BCNT4) );
    zivb U342 ( .A(BCNT4), .Y(n734) );
    zdffqrb BCNT_reg_3 ( .CK(PCICLK), .D(BCNT462_3), .R(HRST_), .Q(BCNT3) );
    zivb U343 ( .A(BCNT3), .Y(n751) );
    zdffqrb BOUNDRY_T_reg ( .CK(PCICLK), .D(BOUNDRY_T425), .R(HRST_), .Q(
        BOUNDRY_T) );
    zivb U344 ( .A(BOUNDRY_T), .Y(n800) );
    zdffrb BTIMER_reg_2 ( .CK(PCICLK), .D(n830), .R(HRST_), .Q(BTIMER_2), .QN(
        n640) );
    zdffrb BTIMER_reg_4 ( .CK(PCICLK), .D(n829), .R(HRST_), .Q(BTIMER_4), .QN(
        n639) );
    znr3b U345 ( .A(n810), .B(n809), .C(SIZEB4), .Y(n593) );
    znr3b U346 ( .A(MBE2_), .B(MBE1_), .C(n798), .Y(n594) );
    zoa21b U347 ( .A(TXREQ), .B(RFREQ_S), .C(n819), .Y(n595) );
    znr2b U348 ( .A(TFGNT), .B(n816), .Y(n596) );
    znr2b U349 ( .A(n818), .B(n797), .Y(n597) );
    znr2b U350 ( .A(MBE3_), .B(MBE2_), .Y(n598) );
    znr3b U351 ( .A(n640), .B(n806), .C(n807), .Y(n599) );
    zan2b U352 ( .A(n600), .B(n783), .Y(n782) );
    zaoi211d U353 ( .A(n816), .B(n805), .C(n769), .D(n620), .Y(n600) );
    zdffrb BCNT_reg_2 ( .CK(PCICLK), .D(BCNT462_2), .R(HRST_), .Q(BCNT2), .QN(
        n627) );
    zdffqrb BCNT_reg_1 ( .CK(PCICLK), .D(BCNT462_1), .R(HRST_), .Q(BCNT1) );
    zivb U354 ( .A(BCNT1), .Y(n810) );
    zdffrb BCNT_reg_5 ( .CK(PCICLK), .D(BCNT462_5), .R(HRST_), .Q(BCNT5), .QN(
        n622) );
    zdffqrb BCNT_reg_0 ( .CK(PCICLK), .D(BCNT462_0), .R(HRST_), .Q(BCNT0) );
    zivb U355 ( .A(BCNT0), .Y(n809) );
    zdffrb BCNT_reg_9 ( .CK(PCICLK), .D(BCNT462_9), .R(HRST_), .Q(BCNT9), .QN(
        n624) );
    zdffqrb BTIMER_reg_0 ( .CK(PCICLK), .D(BTIMER304_0), .R(HRST_), .Q(
        BTIMER_0) );
    zivb U356 ( .A(BTIMER_0), .Y(n807) );
    zdffqrb BCNT_reg_8 ( .CK(PCICLK), .D(BCNT462_8), .R(HRST_), .Q(BCNT8) );
    zivb U357 ( .A(BCNT8), .Y(n634) );
    znr2b U358 ( .A(n641), .B(n640), .Y(n601) );
    znr2b U359 ( .A(n684), .B(n683), .Y(n602) );
    zan2b U360 ( .A(WPR[3]), .B(n700), .Y(n603) );
    zan2b U361 ( .A(n698), .B(n697), .Y(n604) );
    zan2b U362 ( .A(n670), .B(n610), .Y(n605) );
    zan2b U363 ( .A(n675), .B(n676), .Y(n606) );
    zan2b U364 ( .A(n672), .B(n671), .Y(n607) );
    zor2b U365 ( .A(n679), .B(n678), .Y(n608) );
    zor2b U366 ( .A(n679), .B(n650), .Y(n609) );
    zdffqrb BCNT_reg_7 ( .CK(PCICLK), .D(BCNT462_7), .R(HRST_), .Q(BCNT7) );
    zivb U367 ( .A(BCNT6), .Y(n636) );
    zbfb U368 ( .A(n611), .Y(n610) );
    znd2d U369 ( .A(n613), .B(n614), .Y(n611) );
    zivb U370 ( .A(n610), .Y(n708) );
    zor2b U371 ( .A(BCNT7), .B(BCNT6), .Y(n612) );
    zind2b U372 ( .A(n763), .B(n636), .Y(n756) );
    zdffrb BCNT_reg_6 ( .CK(PCICLK), .D(BCNT462_6), .R(HRST_), .Q(BCNT6), .QN(
        n621) );
    znd2b U373 ( .A(n760), .B(n759), .Y(BCNT_NX_0) );
    zivb U374 ( .A(n760), .Y(n743) );
    znd2d U375 ( .A(n646), .B(n616), .Y(n613) );
    zan2d U376 ( .A(n645), .B(n690), .Y(n616) );
    zan2d U377 ( .A(n677), .B(n676), .Y(n617) );
    zan2b U378 ( .A(n602), .B(n652), .Y(n677) );
    znr2d U379 ( .A(n612), .B(n763), .Y(n618) );
    zivb U380 ( .A(n618), .Y(n754) );
    znd4b U381 ( .A(n637), .B(n636), .C(n635), .D(n634), .Y(BCNTBT20) );
    zxo2b U382 ( .A(BTIMER_1), .B(BTIMER_0), .Y(BTIMER290_1) );
    zxo2b U383 ( .A(n640), .B(n641), .Y(BTIMER290_2) );
    zxo2b U384 ( .A(BTIMER_3), .B(n601), .Y(BTIMER290_3) );
    zxo2b U385 ( .A(n639), .B(n638), .Y(BTIMER290_4) );
    znd2d U386 ( .A(n607), .B(WPR[16]), .Y(n663) );
    znd2d U387 ( .A(n676), .B(WPR[18]), .Y(n664) );
    znd2d U388 ( .A(n606), .B(WPR[20]), .Y(n665) );
    znd2d U389 ( .A(n617), .B(n642), .Y(n667) );
    znd2d U390 ( .A(n604), .B(WPR[8]), .Y(n669) );
    znd2d U391 ( .A(n644), .B(n643), .Y(n700) );
    znd2d U392 ( .A(n645), .B(n646), .Y(n643) );
    znd2d U393 ( .A(n702), .B(n740), .Y(n645) );
    znd2d U394 ( .A(n648), .B(n647), .Y(n646) );
    znd2d U395 ( .A(n659), .B(n649), .Y(n647) );
    znd2d U396 ( .A(n703), .B(n741), .Y(n649) );
    znr2d U397 ( .A(n694), .B(n654), .Y(n681) );
    znd4b U398 ( .A(WPR[17]), .B(WPR[16]), .C(WPR[14]), .D(WPR[15]), .Y(n654)
         );
    zan2d U399 ( .A(n782), .B(WPR[0]), .Y(n659) );
    zxo2b U400 ( .A(n720), .B(n660), .Y(WPR_NX_1) );
    zxo2b U401 ( .A(n709), .B(n708), .Y(WPR_NX_10) );
    zxo2b U402 ( .A(WPR[11]), .B(n710), .Y(WPR_NX_11) );
    zxo2b U403 ( .A(n605), .B(WPR[12]), .Y(WPR_NX_12) );
    zxo2b U404 ( .A(n695), .B(n661), .Y(WPR_NX_13) );
    zxo2b U405 ( .A(n689), .B(n674), .Y(WPR_NX_14) );
    zxo2b U406 ( .A(n691), .B(n662), .Y(WPR_NX_15) );
    zxo2b U407 ( .A(n607), .B(WPR[16]), .Y(WPR_NX_16) );
    zxo2b U408 ( .A(n688), .B(n663), .Y(WPR_NX_17) );
    zxo2b U409 ( .A(n686), .B(n682), .Y(WPR_NX_18) );
    zxo2b U410 ( .A(n687), .B(n664), .Y(WPR_NX_19) );
    zxo2b U411 ( .A(n606), .B(WPR[20]), .Y(WPR_NX_20) );
    zxo2b U412 ( .A(n685), .B(n665), .Y(WPR_NX_21) );
    zxo2b U413 ( .A(n711), .B(n726), .Y(WPR_NX_22) );
    zxo2b U414 ( .A(WPR[23]), .B(n712), .Y(WPR_NX_23) );
    zxo2b U415 ( .A(WPR[24]), .B(n727), .Y(WPR_NX_24) );
    zxo2b U416 ( .A(WPR[25]), .B(n714), .Y(WPR_NX_25) );
    zxo2b U417 ( .A(n617), .B(WPR[26]), .Y(WPR_NX_26) );
    zxo2b U418 ( .A(n680), .B(n666), .Y(WPR_NX_27) );
    zxo2b U419 ( .A(WPR[28]), .B(n724), .Y(WPR_NX_28) );
    zxo2b U420 ( .A(n678), .B(n667), .Y(WPR_NX_29) );
    zxo2b U421 ( .A(n721), .B(WPR[30]), .Y(WPR_NX_30) );
    zxo2b U422 ( .A(WPR[31]), .B(n715), .Y(WPR_NX_31) );
    zxo2b U423 ( .A(WPR[4]), .B(n603), .Y(WPR_NX_4) );
    zxo2b U424 ( .A(n701), .B(n668), .Y(WPR_NX_5) );
    zxo2b U425 ( .A(n716), .B(n717), .Y(WPR_NX_6) );
    zxo2b U426 ( .A(WPR[7]), .B(n718), .Y(WPR_NX_7) );
    zxo2b U427 ( .A(n604), .B(WPR[8]), .Y(WPR_NX_8) );
    zxo2b U428 ( .A(n696), .B(n669), .Y(WPR_NX_9) );
    znd2d U429 ( .A(n611), .B(n673), .Y(n674) );
    znd2d U430 ( .A(n676), .B(n602), .Y(n726) );
    znd2d U431 ( .A(n677), .B(n676), .Y(n723) );
    znd2d U432 ( .A(n611), .B(n681), .Y(n682) );
    zxo2b U433 ( .A(n705), .B(n704), .Y(WPR_NX_2) );
    zxo2b U434 ( .A(n707), .B(n706), .Y(WPR_NX_3) );
    znr2d U435 ( .A(n709), .B(n708), .Y(n710) );
    znr2d U436 ( .A(n711), .B(n726), .Y(n712) );
    znr2d U437 ( .A(n726), .B(n713), .Y(n714) );
    znr2d U438 ( .A(n723), .B(n609), .Y(n715) );
    znr2d U439 ( .A(n717), .B(n716), .Y(n718) );
    zinr2b U440 ( .A(n720), .B(n719), .Y(WPR_NX_0) );
    znr2d U441 ( .A(n723), .B(n608), .Y(n721) );
    znr2d U442 ( .A(n723), .B(n722), .Y(n724) );
    znd2d U443 ( .A(n728), .B(n729), .Y(n738) );
    znd2d U444 ( .A(BCNT2), .B(n740), .Y(n733) );
    znd2d U445 ( .A(n731), .B(n730), .Y(n729) );
    znd2d U446 ( .A(n732), .B(n760), .Y(n730) );
    znd2d U447 ( .A(BCNT1), .B(n741), .Y(n731) );
    znd2d U448 ( .A(n782), .B(n809), .Y(n760) );
    zan2d U449 ( .A(n733), .B(n751), .Y(n739) );
    zxo2b U450 ( .A(BCNT10), .B(n747), .Y(BCNT_NX_10) );
    zxo2b U451 ( .A(n624), .B(n758), .Y(BCNT_NX_9) );
    znd2d U452 ( .A(n618), .B(n735), .Y(n758) );
    znd2d U453 ( .A(n737), .B(n736), .Y(n763) );
    znd2d U454 ( .A(n739), .B(n738), .Y(n750) );
    zxo2b U455 ( .A(n744), .B(n743), .Y(BCNT_NX_1) );
    zxo2b U456 ( .A(n746), .B(n745), .Y(BCNT_NX_2) );
    znr2d U457 ( .A(BCNT9), .B(n758), .Y(n747) );
    znr2d U458 ( .A(n749), .B(n748), .Y(n752) );
    zoai21b U459 ( .A(n752), .B(n751), .C(n750), .Y(BCNT_NX_3) );
    znd2d U460 ( .A(n756), .B(n755), .Y(BCNT_NX_6) );
    zoai21b U461 ( .A(n764), .B(n622), .C(n763), .Y(BCNT_NX_5) );
    znd4b U462 ( .A(n768), .B(n767), .C(n766), .D(n765), .Y(SIZEB4) );
    zao21b U463 ( .A(FBE_[2]), .B(n596), .C(n773), .Y(MBE2_) );
    zao222b U464 ( .A(WPR[1]), .B(TFGNT), .C(n774), .D(TFGNT), .E(FBE_[1]), 
        .F(n596), .Y(MBE1_) );
    zoa21d U465 ( .A(NEARBEND), .B(n777), .C(TXFIFO), .Y(TFCOMPL) );
    zoa21d U466 ( .A(n780), .B(n781), .C(n600), .Y(n779) );
    zan4b U467 ( .A(n785), .B(n786), .C(n598), .D(n600), .Y(n784) );
    zao22d U468 ( .A(BUFPTR1[0]), .B(n853), .C(WPR_NX_0), .D(n828), .Y(
        WPR387_0) );
    zao22d U469 ( .A(BUFPTR1[1]), .B(n854), .C(WPR_NX_1), .D(n787), .Y(
        WPR387_1) );
    zao22d U470 ( .A(BUFPTR1[2]), .B(n851), .C(WPR_NX_2), .D(n828), .Y(
        WPR387_2) );
    zao22d U471 ( .A(BUFPTR1[3]), .B(n853), .C(WPR_NX_3), .D(n787), .Y(
        WPR387_3) );
    zao22d U472 ( .A(BUFPTR1[4]), .B(n854), .C(WPR_NX_4), .D(n828), .Y(
        WPR387_4) );
    zao22d U473 ( .A(BUFPTR1[5]), .B(n852), .C(WPR_NX_5), .D(n787), .Y(
        WPR387_5) );
    zao22d U474 ( .A(BUFPTR1[6]), .B(n851), .C(WPR_NX_6), .D(n828), .Y(
        WPR387_6) );
    zao22d U475 ( .A(BUFPTR1[7]), .B(n853), .C(WPR_NX_7), .D(n787), .Y(
        WPR387_7) );
    zao22d U476 ( .A(BUFPTR1[8]), .B(n854), .C(WPR_NX_8), .D(n828), .Y(
        WPR387_8) );
    zao22d U477 ( .A(n853), .B(BUFPTR1[9]), .C(n787), .D(WPR_NX_9), .Y(
        WPR387_9) );
    zao22d U478 ( .A(BUFPTR1[10]), .B(n852), .C(WPR_NX_10), .D(n787), .Y(
        WPR387_10) );
    zao22d U479 ( .A(BUFPTR1[11]), .B(n851), .C(WPR_NX_11), .D(n828), .Y(
        WPR387_11) );
    zao222b U480 ( .A(n831), .B(n788), .C(BUFPTR1[12]), .D(n852), .E(WPR_NX_12
        ), .F(n787), .Y(WPR387_12) );
    zao222b U481 ( .A(n832), .B(n788), .C(BUFPTR1[13]), .D(n853), .E(WPR_NX_13
        ), .F(n828), .Y(WPR387_13) );
    zao222b U482 ( .A(n833), .B(n788), .C(BUFPTR1[14]), .D(n854), .E(WPR_NX_14
        ), .F(n787), .Y(WPR387_14) );
    zao222b U483 ( .A(n834), .B(n788), .C(BUFPTR1[15]), .D(n851), .E(WPR_NX_15
        ), .F(n828), .Y(WPR387_15) );
    zao222b U484 ( .A(n835), .B(n788), .C(BUFPTR1[16]), .D(n852), .E(WPR_NX_16
        ), .F(n787), .Y(WPR387_16) );
    zao222b U485 ( .A(n836), .B(n788), .C(BUFPTR1[17]), .D(n853), .E(WPR_NX_17
        ), .F(n828), .Y(WPR387_17) );
    zao222b U486 ( .A(n837), .B(n788), .C(BUFPTR1[18]), .D(n854), .E(WPR_NX_18
        ), .F(n787), .Y(WPR387_18) );
    zao222b U487 ( .A(n838), .B(n788), .C(BUFPTR1[19]), .D(n851), .E(WPR_NX_19
        ), .F(n828), .Y(WPR387_19) );
    zao222b U488 ( .A(n839), .B(n788), .C(BUFPTR1[20]), .D(n852), .E(WPR_NX_20
        ), .F(n787), .Y(WPR387_20) );
    zao222b U489 ( .A(n840), .B(n788), .C(BUFPTR1[21]), .D(n853), .E(WPR_NX_21
        ), .F(n828), .Y(WPR387_21) );
    zao222b U490 ( .A(n841), .B(n788), .C(BUFPTR1[22]), .D(n854), .E(WPR_NX_22
        ), .F(n787), .Y(WPR387_22) );
    zao222b U491 ( .A(n842), .B(n788), .C(BUFPTR1[23]), .D(n851), .E(WPR_NX_23
        ), .F(n828), .Y(WPR387_23) );
    zao222b U492 ( .A(n843), .B(n788), .C(BUFPTR1[24]), .D(n852), .E(WPR_NX_24
        ), .F(n787), .Y(WPR387_24) );
    zao222b U493 ( .A(n844), .B(n788), .C(BUFPTR1[25]), .D(n853), .E(WPR_NX_25
        ), .F(n828), .Y(WPR387_25) );
    zao222b U494 ( .A(n845), .B(n788), .C(BUFPTR1[26]), .D(n854), .E(WPR_NX_26
        ), .F(n787), .Y(WPR387_26) );
    zao222b U495 ( .A(n846), .B(n788), .C(BUFPTR1[27]), .D(n851), .E(WPR_NX_27
        ), .F(n828), .Y(WPR387_27) );
    zao222b U496 ( .A(n847), .B(n788), .C(BUFPTR1[28]), .D(n852), .E(WPR_NX_28
        ), .F(n787), .Y(WPR387_28) );
    zao222b U497 ( .A(n848), .B(n788), .C(BUFPTR1[29]), .D(n853), .E(WPR_NX_29
        ), .F(n828), .Y(WPR387_29) );
    zao222b U498 ( .A(n849), .B(n788), .C(BUFPTR1[30]), .D(n854), .E(WPR_NX_30
        ), .F(n787), .Y(WPR387_30) );
    zao22d U500 ( .A(n595), .B(BTIMER_3), .C(BTIMER290_3), .D(n789), .Y(
        BTIMER304_3) );
    zao22d U502 ( .A(n595), .B(BTIMER_1), .C(BTIMER290_1), .D(n789), .Y(
        BTIMER304_1) );
    zao22d U503 ( .A(n595), .B(BTIMER_0), .C(n807), .D(n789), .Y(BTIMER304_0)
         );
    zoa21d U504 ( .A(n599), .B(FCFG), .C(BTIMER_3), .Y(n790) );
    zcx7b U505 ( .A(n793), .B(n794), .C(WPR_NX_31), .D(n795), .E(n796), .Y(
        WPR387_31) );
    zxo2b U506 ( .A(MBE2_), .B(n785), .Y(n797) );
    zxo2b U507 ( .A(MBE3_), .B(n785), .Y(n798) );
    zor2d U508 ( .A(n851), .B(BOUNDRY_T), .Y(n799) );
    zor2d U509 ( .A(n852), .B(n800), .Y(n802) );
    zao211b U510 ( .A(FCFG), .B(n599), .C(BTIMER_4), .D(n790), .Y(n777) );
    zor3b U511 ( .A(BCNT1), .B(n809), .C(SIZEB4), .Y(n815) );
    zor3b U512 ( .A(BCNT0), .B(n810), .C(SIZEB4), .Y(n817) );
    znd5d U513 ( .A(DIS_BURST), .B(PMSTR), .C(RFREQ_S), .D(RFGNT), .E(n619), 
        .Y(n819) );
    zxo2b U514 ( .A(n818), .B(n786), .Y(n792) );
    zxo2b U515 ( .A(BTIMER_3), .B(FCFG), .Y(n771) );
    zmux21hd U516 ( .A(n840), .B(BUFPTR2[21]), .S(n852), .Y(BUFPTR2_LT363_9)
         );
    zmux21hd U517 ( .A(n839), .B(BUFPTR2[20]), .S(n853), .Y(BUFPTR2_LT363_8)
         );
    zmux21hd U518 ( .A(n838), .B(BUFPTR2[19]), .S(n854), .Y(BUFPTR2_LT363_7)
         );
    zmux21hd U519 ( .A(n837), .B(BUFPTR2[18]), .S(n852), .Y(BUFPTR2_LT363_6)
         );
    zmux21hd U520 ( .A(n836), .B(BUFPTR2[17]), .S(n853), .Y(BUFPTR2_LT363_5)
         );
    zmux21hd U521 ( .A(n835), .B(BUFPTR2[16]), .S(n854), .Y(BUFPTR2_LT363_4)
         );
    zmux21hd U522 ( .A(n834), .B(BUFPTR2[15]), .S(n851), .Y(BUFPTR2_LT363_3)
         );
    zmux21hd U523 ( .A(n833), .B(BUFPTR2[14]), .S(n852), .Y(BUFPTR2_LT363_2)
         );
    zmux21hd U524 ( .A(n850), .B(BUFPTR2[31]), .S(n853), .Y(BUFPTR2_LT363_19)
         );
    zmux21hd U525 ( .A(n849), .B(BUFPTR2[30]), .S(n854), .Y(BUFPTR2_LT363_18)
         );
    zmux21hd U526 ( .A(n848), .B(BUFPTR2[29]), .S(n851), .Y(BUFPTR2_LT363_17)
         );
    zmux21hd U527 ( .A(n847), .B(BUFPTR2[28]), .S(n852), .Y(BUFPTR2_LT363_16)
         );
    zmux21hd U528 ( .A(n846), .B(BUFPTR2[27]), .S(n853), .Y(BUFPTR2_LT363_15)
         );
    zmux21hd U529 ( .A(n845), .B(BUFPTR2[26]), .S(n854), .Y(BUFPTR2_LT363_14)
         );
    zmux21hd U530 ( .A(n844), .B(BUFPTR2[25]), .S(n851), .Y(BUFPTR2_LT363_13)
         );
    zmux21hd U531 ( .A(n843), .B(BUFPTR2[24]), .S(n852), .Y(BUFPTR2_LT363_12)
         );
    zmux21hd U532 ( .A(n842), .B(BUFPTR2[23]), .S(n853), .Y(BUFPTR2_LT363_11)
         );
    zmux21hd U533 ( .A(n841), .B(BUFPTR2[22]), .S(n854), .Y(BUFPTR2_LT363_10)
         );
    zmux21hd U534 ( .A(n832), .B(BUFPTR2[13]), .S(n851), .Y(BUFPTR2_LT363_1)
         );
    zmux21hd U535 ( .A(n831), .B(BUFPTR2[12]), .S(n852), .Y(BUFPTR2_LT363_0)
         );
    zmux21hd U536 ( .A(BCNT_NX_9), .B(MAXLEN[9]), .S(n853), .Y(BCNT462_9) );
    zmux21hd U537 ( .A(BCNT_NX_8), .B(MAXLEN[8]), .S(n854), .Y(BCNT462_8) );
    zmux21hd U538 ( .A(BCNT_NX_7), .B(MAXLEN[7]), .S(n851), .Y(BCNT462_7) );
    zmux21hd U539 ( .A(BCNT_NX_6), .B(MAXLEN[6]), .S(n852), .Y(BCNT462_6) );
    zmux21hd U540 ( .A(BCNT_NX_5), .B(MAXLEN[5]), .S(n853), .Y(BCNT462_5) );
    zmux21hd U541 ( .A(BCNT_NX_4), .B(MAXLEN[4]), .S(n854), .Y(BCNT462_4) );
    zmux21hd U542 ( .A(BCNT_NX_3), .B(MAXLEN[3]), .S(n851), .Y(BCNT462_3) );
    zmux21hd U543 ( .A(BCNT_NX_2), .B(MAXLEN[2]), .S(n852), .Y(BCNT462_2) );
    zmux21hd U544 ( .A(BCNT_NX_10), .B(MAXLEN[10]), .S(n853), .Y(BCNT462_10)
         );
    zmux21hd U545 ( .A(BCNT_NX_1), .B(MAXLEN[1]), .S(n854), .Y(BCNT462_1) );
    zmux21hd U546 ( .A(BCNT_NX_0), .B(MAXLEN[0]), .S(n851), .Y(BCNT462_0) );
    zan2d U547 ( .A(n824), .B(n799), .Y(n795) );
    zao21b U548 ( .A(n598), .B(MBE0_), .C(n594), .Y(n781) );
    zor6b U549 ( .A(BCNT6), .B(BCNT10), .C(BCNT9), .D(BCNT5), .E(BCNT8), .F(
        BCNT7), .Y(n776) );
    zivf U550 ( .A(n802), .Y(n788) );
    zor2d U551 ( .A(n801), .B(n802), .Y(n796) );
    zivf U552 ( .A(n796), .Y(n794) );
    znd2d U553 ( .A(BUFPTR1[31]), .B(n851), .Y(n824) );
    zivf U554 ( .A(n824), .Y(n793) );
    zoai22b U555 ( .A(WPR[0]), .B(n815), .C(WPR[1]), .D(n821), .Y(n772) );
    zor3b U556 ( .A(n593), .B(SIZEB4), .C(n812), .Y(n827) );
    zao21b U557 ( .A(WPR[0]), .B(n827), .C(WPR[1]), .Y(n775) );
    zao211b U558 ( .A(n597), .B(MBE1_), .C(n594), .D(n791), .Y(n783) );
    zao21b U559 ( .A(n815), .B(n826), .C(n805), .Y(n822) );
    zivl U560 ( .A(n799), .Y(n787) );
    zivl U561 ( .A(n799), .Y(n828) );
    zbfb U562 ( .A(BTIMER304_4), .Y(n829) );
    zao22b U563 ( .A(BTIMER_4), .B(n595), .C(n789), .D(BTIMER290_4), .Y(
        BTIMER304_4) );
    zbfb U564 ( .A(BTIMER304_2), .Y(n830) );
    zao22b U565 ( .A(n595), .B(BTIMER_2), .C(BTIMER290_2), .D(n789), .Y(
        BTIMER304_2) );
    zbfb U566 ( .A(BUFPTR2_LT_0), .Y(n831) );
    zbfb U567 ( .A(BUFPTR2_LT_1), .Y(n832) );
    zbfb U568 ( .A(BUFPTR2_LT_2), .Y(n833) );
    zbfb U569 ( .A(BUFPTR2_LT_3), .Y(n834) );
    zbfb U570 ( .A(BUFPTR2_LT_4), .Y(n835) );
    zbfb U571 ( .A(BUFPTR2_LT_5), .Y(n836) );
    zbfb U572 ( .A(BUFPTR2_LT_6), .Y(n837) );
    zbfb U573 ( .A(BUFPTR2_LT_7), .Y(n838) );
    zbfb U574 ( .A(BUFPTR2_LT_8), .Y(n839) );
    zbfb U575 ( .A(BUFPTR2_LT_9), .Y(n840) );
    zbfb U576 ( .A(BUFPTR2_LT_10), .Y(n841) );
    zbfb U577 ( .A(BUFPTR2_LT_11), .Y(n842) );
    zbfb U578 ( .A(BUFPTR2_LT_12), .Y(n843) );
    zbfb U579 ( .A(BUFPTR2_LT_13), .Y(n844) );
    zbfb U580 ( .A(BUFPTR2_LT_14), .Y(n845) );
    zbfb U581 ( .A(BUFPTR2_LT_15), .Y(n846) );
    zbfb U582 ( .A(BUFPTR2_LT_16), .Y(n847) );
    zbfb U583 ( .A(BUFPTR2_LT_17), .Y(n848) );
    zbfb U584 ( .A(BUFPTR2_LT_18), .Y(n849) );
    zbfb U585 ( .A(BUFPTR2_LT_19), .Y(n850) );
    zbfh U586 ( .A(WPRLD), .Y(n851) );
    zbfh U587 ( .A(WPRLD), .Y(n852) );
    zbfh U588 ( .A(WPRLD), .Y(n853) );
    zbfh U589 ( .A(WPRLD), .Y(n854) );
endmodule


module HS_BMUX ( WPR, FFRDPCI, HCIADR, HCIADD, FIFOGNT, HCIGNT, MA, MWD );
input  [31:0] WPR;
input  [31:0] FFRDPCI;
output [31:0] MA;
input  [31:0] HCIADD;
output [31:0] MWD;
input  [31:0] HCIADR;
input  FIFOGNT, HCIGNT;
    wire n48, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, 
        n63, n64, n65, n66, n67;
    assign MA[1] = 1'b0;
    assign MA[0] = 1'b0;
    zmux21hb U9 ( .A(HCIADR[2]), .B(WPR[2]), .S(n48), .Y(MA[2]) );
    zmux21hb U10 ( .A(HCIADR[3]), .B(WPR[3]), .S(n48), .Y(MA[3]) );
    zymx24hb U11 ( .A1(HCIADR[31]), .A2(HCIADR[30]), .A3(HCIADR[29]), .A4(
        HCIADR[28]), .B1(WPR[31]), .B2(WPR[30]), .B3(WPR[29]), .B4(WPR[28]), 
        .S(n48), .Y1(MA[31]), .Y2(MA[30]), .Y3(MA[29]), .Y4(MA[28]) );
    zymx24hb U12 ( .A1(HCIADR[27]), .A2(HCIADR[26]), .A3(HCIADR[25]), .A4(
        HCIADR[24]), .B1(WPR[27]), .B2(WPR[26]), .B3(WPR[25]), .B4(WPR[24]), 
        .S(n48), .Y1(MA[27]), .Y2(MA[26]), .Y3(MA[25]), .Y4(MA[24]) );
    zymx24hb U13 ( .A1(HCIADR[23]), .A2(HCIADR[22]), .A3(HCIADR[21]), .A4(
        HCIADR[20]), .B1(WPR[23]), .B2(WPR[22]), .B3(WPR[21]), .B4(WPR[20]), 
        .S(n48), .Y1(MA[23]), .Y2(MA[22]), .Y3(MA[21]), .Y4(MA[20]) );
    zymx24hb U14 ( .A1(HCIADR[19]), .A2(HCIADR[18]), .A3(HCIADR[17]), .A4(
        HCIADR[16]), .B1(WPR[19]), .B2(WPR[18]), .B3(WPR[17]), .B4(WPR[16]), 
        .S(n48), .Y1(MA[19]), .Y2(MA[18]), .Y3(MA[17]), .Y4(MA[16]) );
    zymx24hb U15 ( .A1(HCIADR[15]), .A2(HCIADR[14]), .A3(HCIADR[13]), .A4(
        HCIADR[12]), .B1(WPR[15]), .B2(WPR[14]), .B3(WPR[13]), .B4(WPR[12]), 
        .S(n48), .Y1(MA[15]), .Y2(MA[14]), .Y3(MA[13]), .Y4(MA[12]) );
    zymx24hb U16 ( .A1(HCIADR[11]), .A2(HCIADR[10]), .A3(HCIADR[9]), .A4(
        HCIADR[8]), .B1(WPR[11]), .B2(WPR[10]), .B3(WPR[9]), .B4(WPR[8]), .S(
        n48), .Y1(MA[11]), .Y2(MA[10]), .Y3(MA[9]), .Y4(MA[8]) );
    zymx24hb U17 ( .A1(HCIADR[7]), .A2(HCIADR[6]), .A3(HCIADR[5]), .A4(HCIADR
        [4]), .B1(WPR[7]), .B2(WPR[6]), .B3(WPR[5]), .B4(WPR[4]), .S(n48), 
        .Y1(MA[7]), .Y2(MA[6]), .Y3(MA[5]), .Y4(MA[4]) );
    zao22b U18 ( .A(FFRDPCI[0]), .B(FIFOGNT), .C(HCIADD[0]), .D(n66), .Y(MWD
        [0]) );
    zao22b U19 ( .A(FFRDPCI[1]), .B(FIFOGNT), .C(HCIADD[1]), .D(n66), .Y(MWD
        [1]) );
    zao22b U20 ( .A(FFRDPCI[2]), .B(FIFOGNT), .C(HCIADD[2]), .D(n66), .Y(MWD
        [2]) );
    zao21b U21 ( .A(HCIADD[3]), .B(n67), .C(n52), .Y(MWD[3]) );
    zao21b U22 ( .A(FFRDPCI[3]), .B(n48), .C(n51), .Y(n52) );
    zao21b U23 ( .A(HCIADD[4]), .B(n67), .C(n53), .Y(MWD[4]) );
    zao21b U24 ( .A(FFRDPCI[4]), .B(n48), .C(n51), .Y(n53) );
    zao21b U25 ( .A(HCIADD[5]), .B(n66), .C(n54), .Y(MWD[5]) );
    zao21b U26 ( .A(FFRDPCI[5]), .B(n48), .C(n51), .Y(n54) );
    zao21b U27 ( .A(HCIADD[6]), .B(n67), .C(n55), .Y(MWD[6]) );
    zao21b U28 ( .A(FFRDPCI[6]), .B(n48), .C(n51), .Y(n55) );
    zao22b U29 ( .A(FFRDPCI[7]), .B(FIFOGNT), .C(HCIADD[7]), .D(n66), .Y(MWD
        [7]) );
    zao22b U30 ( .A(FFRDPCI[8]), .B(FIFOGNT), .C(HCIADD[8]), .D(n67), .Y(MWD
        [8]) );
    zao21b U31 ( .A(n67), .B(HCIADD[9]), .C(n56), .Y(MWD[9]) );
    zao21b U32 ( .A(HCIADD[10]), .B(n67), .C(n57), .Y(MWD[10]) );
    zao21b U33 ( .A(FFRDPCI[10]), .B(n48), .C(n51), .Y(n57) );
    zao22b U34 ( .A(FFRDPCI[11]), .B(FIFOGNT), .C(HCIADD[11]), .D(n66), .Y(MWD
        [11]) );
    zao21b U35 ( .A(HCIADD[12]), .B(n66), .C(n58), .Y(MWD[12]) );
    zao21b U36 ( .A(FFRDPCI[12]), .B(n48), .C(n51), .Y(n58) );
    zao22b U37 ( .A(FFRDPCI[13]), .B(FIFOGNT), .C(HCIADD[13]), .D(n67), .Y(MWD
        [13]) );
    zao21b U38 ( .A(HCIADD[14]), .B(n67), .C(n59), .Y(MWD[14]) );
    zao21b U39 ( .A(FFRDPCI[14]), .B(n48), .C(n51), .Y(n59) );
    zao22b U40 ( .A(FFRDPCI[15]), .B(FIFOGNT), .C(HCIADD[15]), .D(n67), .Y(MWD
        [15]) );
    zao22b U41 ( .A(FFRDPCI[16]), .B(FIFOGNT), .C(HCIADD[16]), .D(n67), .Y(MWD
        [16]) );
    zao22b U42 ( .A(FFRDPCI[17]), .B(FIFOGNT), .C(HCIADD[17]), .D(n67), .Y(MWD
        [17]) );
    zao21b U43 ( .A(HCIADD[18]), .B(n67), .C(n60), .Y(MWD[18]) );
    zao21b U44 ( .A(FFRDPCI[18]), .B(n48), .C(n51), .Y(n60) );
    zao22b U45 ( .A(FFRDPCI[19]), .B(FIFOGNT), .C(HCIADD[19]), .D(n66), .Y(MWD
        [19]) );
    zao21b U46 ( .A(HCIADD[20]), .B(n67), .C(n61), .Y(MWD[20]) );
    zao21b U47 ( .A(FFRDPCI[20]), .B(n48), .C(n51), .Y(n61) );
    zao21b U48 ( .A(HCIADD[21]), .B(n67), .C(n62), .Y(MWD[21]) );
    zao21b U49 ( .A(FFRDPCI[21]), .B(FIFOGNT), .C(n51), .Y(n62) );
    zao22b U50 ( .A(FFRDPCI[22]), .B(FIFOGNT), .C(HCIADD[22]), .D(n66), .Y(MWD
        [22]) );
    zao22b U51 ( .A(FFRDPCI[23]), .B(FIFOGNT), .C(HCIADD[23]), .D(n66), .Y(MWD
        [23]) );
    zao22b U52 ( .A(FFRDPCI[24]), .B(FIFOGNT), .C(HCIADD[24]), .D(n66), .Y(MWD
        [24]) );
    zao21b U53 ( .A(HCIADD[25]), .B(n67), .C(n63), .Y(MWD[25]) );
    zao21b U54 ( .A(FFRDPCI[25]), .B(n48), .C(n51), .Y(n63) );
    zao22b U55 ( .A(FFRDPCI[26]), .B(FIFOGNT), .C(HCIADD[26]), .D(n66), .Y(MWD
        [26]) );
    zao22b U56 ( .A(FFRDPCI[27]), .B(FIFOGNT), .C(HCIADD[27]), .D(n66), .Y(MWD
        [27]) );
    zao21b U57 ( .A(HCIADD[28]), .B(n67), .C(n64), .Y(MWD[28]) );
    zao21b U58 ( .A(FFRDPCI[28]), .B(n48), .C(n51), .Y(n64) );
    zao22b U59 ( .A(FFRDPCI[29]), .B(FIFOGNT), .C(HCIADD[29]), .D(n66), .Y(MWD
        [29]) );
    zao22b U60 ( .A(FFRDPCI[30]), .B(FIFOGNT), .C(HCIADD[30]), .D(n66), .Y(MWD
        [30]) );
    zao22b U61 ( .A(FFRDPCI[31]), .B(FIFOGNT), .C(HCIADD[31]), .D(n66), .Y(MWD
        [31]) );
    zivb U62 ( .A(HCIGNT), .Y(n65) );
    zbfb U63 ( .A(n50), .Y(n67) );
    zbfb U64 ( .A(n50), .Y(n66) );
    znr2b U65 ( .A(FIFOGNT), .B(n65), .Y(n50) );
    znr2b U66 ( .A(FIFOGNT), .B(HCIGNT), .Y(n51) );
    zbfb U67 ( .A(FIFOGNT), .Y(n48) );
    zao21b U68 ( .A(FIFOGNT), .B(FFRDPCI[9]), .C(n51), .Y(n56) );
endmodule


module HS_BMUIF ( CREQ, MRDY_, CACHEN, COMPL, MSWR, MRDMPLZ, XMITNULL, WPRLD, 
    PCIREAD, PCIWRT, NEARFEMP, NEARFULL, TXTHRESH, RXTHRESH, MYPMACK, WPR1, 
    WPR0, BCNTBT40, MAXLEN, CACHLN7, CACHLN6, CACHLN5, CACHLN4, CACHLN3, 
    CACHLN2, CACHLN1, CACHLN0, CAHCFG_, RFCOMPL, TFCOMPL, BUFEND, HCIGNT, 
    FIFOGNT, FEMPTY, FCOUNT, XMITSTRT, RXSTRT, TFGNT, RFGNT, TXREQ, RXREQ, 
    RFREQ_S, FCFG, MWRMEN, HCIREQ, HCICOMPL, HCIMWR, HCIMRDY, PMSTR, MADDR, 
    PCI1WAIT, TXFIFO, RXFIFO, EOTQ, RDYACK, PCICLK, HRST_, TADOE, UADOE_, 
    BOUNDRY, BOUNDRY_T, DIS_BURST, ZEROLEN, FIFO_OK );
input  [10:0] MAXLEN;
input  [8:0] FCOUNT;
input  WPR1, WPR0, BCNTBT40, CACHLN7, CACHLN6, CACHLN5, CACHLN4, CACHLN3, 
    CACHLN2, CACHLN1, CACHLN0, CAHCFG_, RFCOMPL, TFCOMPL, BUFEND, HCIGNT, 
    FIFOGNT, FEMPTY, XMITSTRT, RXSTRT, TFGNT, RFGNT, TXREQ, RXREQ, RFREQ_S, 
    FCFG, MWRMEN, HCIREQ, HCICOMPL, HCIMWR, HCIMRDY, PMSTR, MADDR, PCI1WAIT, 
    TXFIFO, RXFIFO, EOTQ, RDYACK, PCICLK, HRST_, TADOE, BOUNDRY, BOUNDRY_T, 
    DIS_BURST, FIFO_OK;
output CREQ, MRDY_, CACHEN, COMPL, MSWR, MRDMPLZ, XMITNULL, WPRLD, PCIREAD, 
    PCIWRT, NEARFEMP, NEARFULL, TXTHRESH, RXTHRESH, MYPMACK, UADOE_, ZEROLEN;
    wire SPAREO6, UP_MARK_4, CREQTURN489, SPAREO0_, UP_MARK_3, SPAREO8, n_36, 
        SPAREO1, SPAREO9, COMPLQ452, SPAREO0, n386, FNOTRDY415, SPAREO7, 
        CREQTURN, SPAREO5, n396, SPAREO2, COMPLQ, SPAREO3, SPAREO1_, UP_MARK_8, 
        n_33, SPAREO4, FNOTRDY, n522, n523, n524, n525, n526, n527, n528, n529, 
        n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
        n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, 
        n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, 
        n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, 
        n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;
    zivb SPARE707 ( .A(SPAREO4), .Y(SPAREO5) );
    zdffrb SPARE700 ( .CK(PCICLK), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE709 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE701 ( .CK(PCICLK), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE708 ( .A(SPAREO5), .Y(SPAREO6) );
    znr3b SPARE706 ( .A(SPAREO2), .B(TXTHRESH), .C(SPAREO0_), .Y(SPAREO4) );
    zoai21b SPARE704 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE703 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zaoi211b SPARE702 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE705 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    znd2b U62 ( .A(n552), .B(n546), .Y(n545) );
    znr2b U63 ( .A(FCOUNT[1]), .B(FCOUNT[2]), .Y(n552) );
    znd2b U64 ( .A(FCOUNT[0]), .B(UP_MARK_8), .Y(n546) );
    znd2b U65 ( .A(UP_MARK_3), .B(n560), .Y(n544) );
    znd2b U66 ( .A(n543), .B(n555), .Y(n542) );
    znd3b U67 ( .A(n550), .B(n549), .C(n548), .Y(n551) );
    znd2b U68 ( .A(n557), .B(n556), .Y(n558) );
    znd2b U69 ( .A(n544), .B(n545), .Y(n557) );
    znd2b U70 ( .A(FCOUNT[3]), .B(n559), .Y(n556) );
    zivb U71 ( .A(n558), .Y(n543) );
    znd3b U72 ( .A(n531), .B(n533), .C(RXFIFO), .Y(n530) );
    zivb U73 ( .A(FCOUNT[1]), .Y(n531) );
    znr2b U74 ( .A(FCOUNT[0]), .B(FCOUNT[2]), .Y(n533) );
    znd2b U75 ( .A(UP_MARK_3), .B(n560), .Y(n529) );
    znd2b U76 ( .A(n554), .B(n553), .Y(n561) );
    zaoi21b U77 ( .A(FCOUNT[4]), .B(n558), .C(n551), .Y(n554) );
    znd2b U78 ( .A(n542), .B(n547), .Y(n553) );
    zan2b U79 ( .A(RXFIFO), .B(n573), .Y(UP_MARK_4) );
    zivb U80 ( .A(FCFG), .Y(n573) );
    zivb U81 ( .A(UP_MARK_4), .Y(n547) );
    znd3b U82 ( .A(n550), .B(n549), .C(n548), .Y(n532) );
    znd2b U83 ( .A(n536), .B(n535), .Y(n537) );
    znd2b U84 ( .A(n529), .B(n530), .Y(n536) );
    znd2b U85 ( .A(FCOUNT[3]), .B(n559), .Y(n535) );
    znr2b U86 ( .A(FCOUNT[8]), .B(n561), .Y(n563) );
    znd2b U87 ( .A(FCOUNT[8]), .B(n561), .Y(n562) );
    znd2b U88 ( .A(n523), .B(n524), .Y(n527) );
    znr2b U89 ( .A(FCOUNT[6]), .B(FCOUNT[2]), .Y(n523) );
    znr2b U90 ( .A(FCOUNT[1]), .B(FCOUNT[0]), .Y(n524) );
    znd2b U91 ( .A(n525), .B(n526), .Y(n528) );
    znr2b U92 ( .A(FCOUNT[4]), .B(FCOUNT[5]), .Y(n525) );
    znr2b U93 ( .A(FCOUNT[7]), .B(FCOUNT[3]), .Y(n526) );
    znd2b U94 ( .A(n534), .B(n522), .Y(n538) );
    zaoi21b U95 ( .A(FCOUNT[4]), .B(n537), .C(n532), .Y(n534) );
    zivb U96 ( .A(n537), .Y(n539) );
    znd2b U97 ( .A(FIFO_OK), .B(RXREQ), .Y(n588) );
    zor2b U98 ( .A(BUFEND), .B(n577), .Y(n589) );
    zivb U99 ( .A(TFGNT), .Y(n577) );
    zan2b U100 ( .A(CREQ), .B(COMPL), .Y(COMPLQ452) );
    zivb U101 ( .A(TADOE), .Y(UADOE_) );
    zan3b U102 ( .A(DIS_BURST), .B(RXFIFO), .C(n572), .Y(RXTHRESH) );
    zan2b U103 ( .A(n386), .B(TXFIFO), .Y(TXTHRESH) );
    znr2b U104 ( .A(FCOUNT[8]), .B(n538), .Y(n541) );
    znd2b U105 ( .A(FCOUNT[8]), .B(n538), .Y(n540) );
    znr8b U106 ( .A(FCOUNT[7]), .B(FCOUNT[3]), .C(FCOUNT[1]), .D(FCOUNT[2]), 
        .E(FCOUNT[6]), .F(FCOUNT[8]), .G(FCOUNT[4]), .H(FCOUNT[5]), .Y(
        NEARFEMP) );
    zor2b U107 ( .A(XMITSTRT), .B(RXSTRT), .Y(WPRLD) );
    zan2b U108 ( .A(TXFIFO), .B(ZEROLEN), .Y(XMITNULL) );
    zivb U109 ( .A(BCNTBT40), .Y(n582) );
    zao22b U110 ( .A(HCIMWR), .B(HCIGNT), .C(FIFOGNT), .D(RXFIFO), .Y(MSWR) );
    zan2b U111 ( .A(TFCOMPL), .B(TFGNT), .Y(n564) );
    zan3b U112 ( .A(n569), .B(n570), .C(n571), .Y(CACHEN) );
    zao33b U113 ( .A(MWRMEN), .B(RFREQ_S), .C(RXFIFO), .D(BCNTBT40), .E(TXREQ), 
        .F(TXFIFO), .Y(n569) );
    zivb U114 ( .A(CAHCFG_), .Y(n570) );
    zivb U115 ( .A(n568), .Y(n571) );
    zmux21lb U116 ( .A(n586), .B(n587), .S(FIFOGNT), .Y(MRDY_) );
    zor2b U117 ( .A(HCIMRDY), .B(n578), .Y(n586) );
    zivb U118 ( .A(HCIGNT), .Y(n578) );
    zivb U119 ( .A(HCIMRDY), .Y(n580) );
    zivb U120 ( .A(TXFIFO), .Y(n566) );
    zivb U121 ( .A(TXREQ), .Y(n583) );
    zivb U122 ( .A(RFGNT), .Y(n576) );
    zdffqrb CREQTURN_reg ( .CK(PCICLK), .D(CREQTURN489), .R(HRST_), .Q(
        CREQTURN) );
    zdffqrb COMPLQ_reg ( .CK(PCICLK), .D(COMPLQ452), .R(HRST_), .Q(COMPLQ) );
    zdffqrb FNOTRDY_reg ( .CK(PCICLK), .D(FNOTRDY415), .R(HRST_), .Q(FNOTRDY)
         );
    zaoi211b U123 ( .A(n584), .B(n585), .C(BOUNDRY_T), .D(CREQTURN), .Y(CREQ)
         );
    znr6b U124 ( .A(MAXLEN[2]), .B(MAXLEN[5]), .C(MAXLEN[6]), .D(MAXLEN[1]), 
        .E(MAXLEN[4]), .F(n579), .Y(ZEROLEN) );
    zivb U125 ( .A(FCOUNT[3]), .Y(n560) );
    zan2b U126 ( .A(FCFG), .B(RXFIFO), .Y(UP_MARK_3) );
    zivb U127 ( .A(UP_MARK_3), .Y(n559) );
    zivb U128 ( .A(FCOUNT[4]), .Y(n555) );
    zivb U129 ( .A(FCOUNT[7]), .Y(n549) );
    zivb U130 ( .A(RXFIFO), .Y(UP_MARK_8) );
    zivb U131 ( .A(FCOUNT[5]), .Y(n550) );
    zivb U132 ( .A(FCOUNT[6]), .Y(n548) );
    zao21b U133 ( .A(n539), .B(n555), .C(UP_MARK_4), .Y(n522) );
    zoai21b U134 ( .A(n528), .B(n527), .C(FCOUNT[8]), .Y(n386) );
    zoai21b U135 ( .A(UP_MARK_8), .B(n541), .C(n540), .Y(NEARFULL) );
    zoai21b U136 ( .A(UP_MARK_8), .B(n563), .C(n562), .Y(n396) );
    zao211b U137 ( .A(HCIGNT), .B(HCICOMPL), .C(n564), .D(n565), .Y(COMPL) );
    zor4b U138 ( .A(CAHCFG_), .B(n566), .C(n567), .D(n568), .Y(MRDMPLZ) );
    zoa211b U139 ( .A(RDYACK), .B(MADDR), .C(PCI1WAIT), .D(FIFOGNT), .Y(
        FNOTRDY415) );
    zoa21d U140 ( .A(RFGNT), .B(TFGNT), .C(BOUNDRY), .Y(n574) );
    zxn2b U141 ( .A(CACHLN3), .B(CACHLN2), .Y(n575) );
    zor6b U142 ( .A(CACHLN4), .B(WPR1), .C(CACHLN6), .D(CACHLN5), .E(CACHLN0), 
        .F(n581), .Y(n568) );
    zao211b U143 ( .A(RFCOMPL), .B(RFGNT), .C(COMPLQ), .D(n574), .Y(n565) );
    zor6b U144 ( .A(MAXLEN[9]), .B(MAXLEN[8]), .C(MAXLEN[3]), .D(MAXLEN[7]), 
        .E(MAXLEN[10]), .F(MAXLEN[0]), .Y(n579) );
    zor4b U145 ( .A(CACHLN7), .B(n575), .C(WPR0), .D(CACHLN1), .Y(n581) );
    zao211b U146 ( .A(DIS_BURST), .B(FCFG), .C(n583), .D(n582), .Y(n567) );
    zcx7b U147 ( .A(n566), .B(n583), .C(n589), .D(HCIREQ), .E(HCIGNT), .Y(n584
        ) );
    zao21b U148 ( .A(NEARFULL), .B(EOTQ), .C(n396), .Y(n572) );
    zor4b U149 ( .A(FEMPTY), .B(n576), .C(UP_MARK_8), .D(n588), .Y(n585) );
    zoai21b U150 ( .A(n578), .B(n580), .C(FNOTRDY), .Y(n587) );
    zan2d S_27 ( .A(RDYACK), .B(TFGNT), .Y(n_36) );
    zan2d S_28 ( .A(n_36), .B(PMSTR), .Y(PCIWRT) );
    zan2d S_115 ( .A(COMPL), .B(RDYACK), .Y(CREQTURN489) );
    zan2d S_26 ( .A(RDYACK), .B(PMSTR), .Y(MYPMACK) );
    zan2d S_24 ( .A(RDYACK), .B(RFGNT), .Y(n_33) );
    zan2d S_25 ( .A(n_33), .B(PMSTR), .Y(PCIREAD) );
endmodule

//	@(#)bmuc.src	1.3	17 May 1997
/******************************************************************
- iterface and data MUX between PCIM engine and data buffer control and UHCI control
Timing Issues:
Design Notes:
	- CACHE : on what case .. assert MRDL MRDM command ??

= HCIADD HCIGNT and data select and be select to MUX to PCI I/F
	- take care of MADOE + TADOE .... drivibility ??

(*) exact dword count in databuf = FCOUNT+1

== I/F from HCI control
1. HCIGNT : Internal arbiter grant DESC DMA
2. DESC : DESC DMA DATA
4. FIFOGNT : Internal arbiter grant FIFO DATADMA
5. HCICOMPL : DESC DMA look ahead complete
6. HCIMWR : DESC DMA WRITE
1. WPR is used by test mode and normal mode

- MRDY_ ???
- HCIMRDY
- diffewrence between HCIREQ and HCICREQ ?? 

*******************************************************************/

module HS_BMUC ( 
		/* output */
		//UAD31O, UAD30O, UAD29O, UAD28O, UAD27O, UAD26O,
                //UAD25O, UAD24O, UAD23O, UAD22O, UAD21O, UAD20O,
                //UAD19O, UAD18O, UAD17O, UAD16O, UAD15O, UAD14O,
                //UAD13O, UAD12O, UAD11O, UAD10O, UAD9O,  UAD8O,
                //UAD7O,  UAD6O,  UAD5O,  UAD4O,  UAD3O,  UAD2O,
                //UAD1O,  UAD0O, 
		MA, MWD,
		/*WPR31, WPR30, WPR29, WPR28, WPR27, WPR26,
                WPR25, WPR24, WPR23, WPR22, WPR21, WPR20,
                WPR19, WPR18, WPR17, WPR16, WPR15, WPR14,
                WPR13, WPR12, WPR11, WPR10, WPR9,  WPR8,
                WPR7,  WPR6,  WPR5,  WPR4,  WPR3,  WPR2,*/
                WPR,
		//BCNT10, BCNT9,  BCNT8, BCNT7,  BCNT6,  BCNT5,  
		//BCNT4,  BCNT3,  BCNT2, BCNT1,  BCNT0,
		MBE3_, MBE2_, MBE1_,MBE0_, CREQ, MRDY_, CACHEN, 
		COMPL, MSWR, MRDMPLZ, XMITNULL, 
		UMORE, UMORE2LN,
		PCIREAD, PCIWRT, HCIGNT, RDMAEND, TDMAEND, 
		//TXTHRESH2,	// added by Chris Lai, 5/5/1999
		TXTHRESH,

		/* input */
		//PSADO31, PSADO30, PSADO29, PSADO28, PSADO27, PSADO26,
                //PSADO25, PSADO24, PSADO23, PSADO22, PSADO21, PSADO20,
                //PSADO19, PSADO18, PSADO17, PSADO16, PSADO15, PSADO14,
                //PSADO13, PSADO12, PSADO11, PSADO10, PSADO9,  PSADO8,
                //PSADO7,  PSADO6,  PSADO5,  PSADO4,  PSADO3,  PSADO2,
                //PSADO1,  PSADO0,

		/*FFDOUT31, FFDOUT30, FFDOUT29, FFDOUT28, FFDOUT27, FFDOUT26,
                FFDOUT25, FFDOUT24, FFDOUT23, FFDOUT22, FFDOUT21, FFDOUT20,
                FFDOUT19, FFDOUT18, FFDOUT17, FFDOUT16, FFDOUT15, FFDOUT14,
                FFDOUT13, FFDOUT12, FFDOUT11, FFDOUT10, FFDOUT9,  FFDOUT8,
                FFDOUT7,  FFDOUT6,  FFDOUT5,  FFDOUT4,  FFDOUT3,  FFDOUT2,
                FFDOUT1,  FFDOUT0, */
		FFRDPCI,

		/*BUFPTR31, BUFPTR30, BUFPTR29, BUFPTR28, BUFPTR27, BUFPTR26,
                BUFPTR25, BUFPTR24, BUFPTR23, BUFPTR22, BUFPTR21, BUFPTR20,
                BUFPTR19, BUFPTR18, BUFPTR17, BUFPTR16, BUFPTR15, BUFPTR14,
                BUFPTR13, BUFPTR12, BUFPTR11, BUFPTR10, BUFPTR9,  BUFPTR8,
                BUFPTR7,  BUFPTR6,  BUFPTR5,  BUFPTR4,  BUFPTR3,  BUFPTR2,
                BUFPTR1,  BUFPTR0,*/
		BUFPTR1, BUFPTR2,

		/*HCIADR31, HCIADR30, HCIADR29, HCIADR28, HCIADR27, HCIADR26,
                HCIADR25, HCIADR24, HCIADR23, HCIADR22, HCIADR21, HCIADR20,
                HCIADR19, HCIADR18, HCIADR17, HCIADR16, HCIADR15, HCIADR14,
                HCIADR13, HCIADR12, HCIADR11, HCIADR10, HCIADR9,  HCIADR8,
                HCIADR7,  HCIADR6,  HCIADR5,  HCIADR4,  HCIADR3,  HCIADR2,
                HCIADR1,  HCIADR0,*/
		HCIADR,
		/*HCIADD31, HCIADD30, HCIADD29, HCIADD28, HCIADD27, HCIADD26,
                HCIADD25, HCIADD24, HCIADD23, HCIADD22, HCIADD21, HCIADD20,
                HCIADD19, HCIADD18, HCIADD17, HCIADD16, HCIADD15, HCIADD14,
                HCIADD13, HCIADD12, HCIADD11, HCIADD10, HCIADD9,  HCIADD8,
                HCIADD7,  HCIADD6,  HCIADD5,  HCIADD4,  HCIADD3,  HCIADD2,
                HCIADD1,  HCIADD0,*/
		HCIADD,
		/*MAXLEN10, MAXLEN9,  MAXLEN8, MAXLEN7,  MAXLEN6,  MAXLEN5,  
		MAXLEN4,  MAXLEN3,  MAXLEN2, MAXLEN1,  MAXLEN0,*/
		MAXLEN,
		CACHLN7,  CACHLN6,  CACHLN5,  CACHLN4,  CACHLN3,  CACHLN2,
                CACHLN1,  CACHLN0, CAHCFG_,

		//FBE3_, FBE2_, FBE1_,FBE0_, 
		FBE_,
		RXPKTEND, FEMPTY, //FCOUNT4,FCOUNT3,FCOUNT2,FCOUNT1,FCOUNT0, 
		FCOUNT,
		QRXERR, MABORTS, TABORTR, XMITSTRT, RXSTRT,
		BUSFREE , UGNTI_,
		/*PMDSEL,*/ MWRMEN, 
		HCIREQ, HCICOMPL, HCIMWR, PMSTR, MADDR, PCI1WAIT, 
		EOTQ, TXFIFO, RXFIFO, RDYACK, //UCBE3O_, UCBE2O_, UCBE1O_,UCBE0O_, 
		FCFG, HCIMRDY, 
		//PCICLK, PCICLK2, HRST_ 
		PCICLK, HRST_,
		DISTXDLY, EOF, 		// by Chris Lai, 6/25/1999
		DISTXDLY2, BMUSM_RST_EN, DBUFERR, DISPFIFO,
		DISRXZERO, BUI_GO, DISPFIFO2,
		ENBMUSMRST,		// by Chris Lai, 10/26/1999
		TADOE, /*MADOE,*/ UADOE_, BOUNDRY, DIS_BURST, FIFO_OK,
		DMA_IDLE, ATPG_ENI
		);

// FIFOACK must be more qualified !!

input		FIFO_OK;
output		UMORE, UMORE2LN;
output		DMA_IDLE;
//input		TEST_PACKET;	// in Test_Packet test mode, BMUC deactivated
output [31:0]   MA, MWD;

input		TADOE, /*MADOE,*/ DIS_BURST;
output		UADOE_, BOUNDRY;
input		DISTXDLY2, BMUSM_RST_EN, DBUFERR, DISPFIFO,
		DISRXZERO, BUI_GO, DISPFIFO2,
		ENBMUSMRST;             // by Chris Lai, 10/26/1999
input		DISTXDLY, EOF;		// by Chris Lai, 6/25/1999
//output		TXTHRESH2;	// added by Chris Lai, 5/5/1999
output		TXTHRESH;	// added by Chris Lai, 5/5/1999
/*
output		UAD31O;
output		UAD30O;
output		UAD29O;
output		UAD28O;
output		UAD27O;
output		UAD26O;

output		UAD25O;
output		UAD24O;
output		UAD23O;
output		UAD22O;
output		UAD21O;
output		UAD20O;

output		UAD19O;
output		UAD18O;
output		UAD17O;
output		UAD16O;
output		UAD15O;
output		UAD14O;

output		UAD13O;
output		UAD12O;
output		UAD11O;
output		UAD10O;
output		UAD9O;
output		UAD8O;

output		UAD7O;
output		UAD6O;
output		UAD5O;
output		UAD4O;
output		UAD3O;
output		UAD2O;

output		UAD1O;
output		UAD0O;

output		WPR31;
output		WPR30;
output		WPR29;
output		WPR28;
output		WPR27;
output		WPR26;

output		WPR25;
output		WPR24;
output		WPR23;
output		WPR22;
output		WPR21;
output		WPR20;

output		WPR19;
output		WPR18;
output		WPR17;
output		WPR16;
output		WPR15;
output		WPR14;

output		WPR13;
output		WPR12;
output		WPR11;
output		WPR10;
output		WPR9;
output		WPR8;

output		WPR7;
output		WPR6;
output		WPR5;
output		WPR4;
output		WPR3;
output		WPR2;

output		WPR1;
output		WPR0;*/
output	[31:0]	WPR;

/*output		BCNT10;
output		BCNT9;
output		BCNT8;
output		BCNT7;
output		BCNT6;
output		BCNT5;

output		BCNT4;
output		BCNT3;
output		BCNT2;
output		BCNT1;
output		BCNT0;*/

output		MBE3_;
output		MBE2_;
output		MBE1_;
output		MBE0_;
output		CREQ;
output		MRDY_;
output		CACHEN;

output		COMPL;
output		MSWR;
output		MRDMPLZ;
output		XMITNULL;

output		PCIREAD;
output		PCIWRT;
output		HCIGNT;
output		RDMAEND;
output		TDMAEND;
/*
input		PSADO31;
input		PSADO30;
input		PSADO29;
input		PSADO28;
input		PSADO27;
input		PSADO26;

input		PSADO25;
input		PSADO24;
input		PSADO23;
input		PSADO22;
input		PSADO21;
input		PSADO20;

input		PSADO19;
input		PSADO18;
input		PSADO17;
input		PSADO16;
input		PSADO15;
input		PSADO14;

input		PSADO13;
input		PSADO12;
input		PSADO11;
input		PSADO10;
input		PSADO9;
input		PSADO8;

input		PSADO7;
input		PSADO6;
input		PSADO5;
input		PSADO4;
input		PSADO3;
input		PSADO2;

input		PSADO1;
input		PSADO0;

input		FFDOUT31;
input		FFDOUT30;
input		FFDOUT29;
input		FFDOUT28;
input		FFDOUT27;
input		FFDOUT26;

input		FFDOUT25;
input		FFDOUT24;
input		FFDOUT23;
input		FFDOUT22;
input		FFDOUT21;
input		FFDOUT20;

input		FFDOUT19;
input		FFDOUT18;
input		FFDOUT17;
input		FFDOUT16;
input		FFDOUT15;
input		FFDOUT14;

input		FFDOUT13;
input		FFDOUT12;
input		FFDOUT11;
input		FFDOUT10;
input		FFDOUT9;
input		FFDOUT8;

input		FFDOUT7;
input		FFDOUT6;
input		FFDOUT5;
input		FFDOUT4;
input		FFDOUT3;
input		FFDOUT2;

input		FFDOUT1;
input		FFDOUT0;*/
input	[31:0]	FFRDPCI;

/*input		BUFPTR31;
input		BUFPTR30;
input		BUFPTR29;
input		BUFPTR28;
input		BUFPTR27;
input		BUFPTR26;

input		BUFPTR25;
input		BUFPTR24;
input		BUFPTR23;
input		BUFPTR22;
input		BUFPTR21;
input		BUFPTR20;

input		BUFPTR19;
input		BUFPTR18;
input		BUFPTR17;
input		BUFPTR16;
input		BUFPTR15;
input		BUFPTR14;

input		BUFPTR13;
input		BUFPTR12;
input		BUFPTR11;
input		BUFPTR10;
input		BUFPTR9;
input		BUFPTR8;

input		BUFPTR7;
input		BUFPTR6;
input		BUFPTR5;
input		BUFPTR4;
input		BUFPTR3;
input		BUFPTR2;

input		BUFPTR1;
input		BUFPTR0;*/
input	[31:0]	BUFPTR1, BUFPTR2;

/*input		HCIADR31;
input		HCIADR30;
input		HCIADR29;
input		HCIADR28;
input		HCIADR27;
input		HCIADR26;

input		HCIADR25;
input		HCIADR24;
input		HCIADR23;
input		HCIADR22;
input		HCIADR21;
input		HCIADR20;

input		HCIADR19;
input		HCIADR18;
input		HCIADR17;
input		HCIADR16;
input		HCIADR15;
input		HCIADR14;

input		HCIADR13;
input		HCIADR12;
input		HCIADR11;
input		HCIADR10;
input		HCIADR9;
input		HCIADR8;

input		HCIADR7;
input		HCIADR6;
input		HCIADR5;
input		HCIADR4;
input		HCIADR3;
input		HCIADR2;

input		HCIADR1;
input		HCIADR0;

input		HCIADD31;
input		HCIADD30;
input		HCIADD29;
input		HCIADD28;
input		HCIADD27;
input		HCIADD26;

input		HCIADD25;
input		HCIADD24;
input		HCIADD23;
input		HCIADD22;
input		HCIADD21;
input		HCIADD20;

input		HCIADD19;
input		HCIADD18;
input		HCIADD17;
input		HCIADD16;
input		HCIADD15;
input		HCIADD14;

input		HCIADD13;
input		HCIADD12;
input		HCIADD11;
input		HCIADD10;
input		HCIADD9;
input		HCIADD8;

input		HCIADD7;
input		HCIADD6;
input		HCIADD5;
input		HCIADD4;
input		HCIADD3;
input		HCIADD2;

input		HCIADD1;
input		HCIADD0;*/
input	[31:0]	HCIADR, HCIADD;

/*input		MAXLEN10;
input		MAXLEN9;
input		MAXLEN8;
input		MAXLEN7;
input		MAXLEN6;
input		MAXLEN5;

input		MAXLEN4;
input		MAXLEN3;
input		MAXLEN2;
input		MAXLEN1;
input		MAXLEN0;*/
input	[10:0]	MAXLEN;

input		CACHLN7;
input		CACHLN6;
input		CACHLN5;
input		CACHLN4;
input		CACHLN3;
input		CACHLN2;

input		CACHLN1;
input		CACHLN0;
input		CAHCFG_;


/*input		FBE3_;
input		FBE2_;
input		FBE1_;
input		FBE0_;*/
input	[3:0]	FBE_;

input		RXPKTEND;
input		FEMPTY;
/*input		FCOUNT4;
input		FCOUNT3;
input		FCOUNT2;
input		FCOUNT1;
input		FCOUNT0;*/
input	[8:0]	FCOUNT;

input		QRXERR;
input		MABORTS;
input		TABORTR;
input		XMITSTRT;
input		RXSTRT;

input		BUSFREE;
input		UGNTI_;

//input		PMDSEL;
input		MWRMEN;

input		HCIREQ;
input		HCICOMPL;
input		HCIMWR;
input		PMSTR;
input		MADDR;
input		PCI1WAIT;

input		EOTQ;
input		TXFIFO;
input		RXFIFO;
input		RDYACK;
//input		UCBE3O_;
//input		UCBE2O_;
//input		UCBE1O_;
//input		UCBE0O_;

input		FCFG;
input		HCIMRDY;

//input		PCICLK, PCICLK2;
input		PCICLK;
input		HRST_;
input		ATPG_ENI;

// wire BMURST_ = HRST_ & ~TEST_PACKET;
//sivb DNT0 ( .A(TEST_PACKET), .Y(TEST_PACKET_) );
//san2b DNT1 ( .A(HRST_), .B(TEST_PACKET_), .Y(BMURST_) );

// #define HRST_ BMURST_





HS_BMUSM HS_BMUSM ( 
		/* output */
		HCIGNT, FIFOGNT, RDMAEND, TDMAEND, TXREQ, RXREQ,
		RFREQ_S, RFLUSH_S,

		/* input */
		EOTQ, XMITSTRT, TXTHRESH, XMITNULL, BUFEND,MABORTS, TABORTR,  
		BUSTMOUT, FEMPTY, MYPMACK,
		RXSTRT, QRXERR, RXTHRESH, RXPKTEND, 
		BUSFREE , 1'b0, HCIREQ,
		PCICLK, HRST_,
		DISTXDLY, EOF,		// by Chris Lai, 6/25/1999
		DISTXDLY2, BMUSM_RST_EN,// by Chris Lai, 10/7/1999
		DBUFERR, DISPFIFO,	// by Chris Lai, 10/6/1999
		ZEROLEN, DISRXZERO,	// by Chris Lai, 10/6/1999
		BUI_GO,			// by Chris Lai, 10/8/1999
		DISPFIFO2, ENBMUSMRST,	// by Chris Lai, 10/18/1999, 69B
		DMA_IDLE, ATPG_ENI,
		FIFO_OK 		// by Chris Lai, 3/18/2003, 104B5
		);


HS_BMUTM HS_BMUTM ( 
		/* output */
		/*WPR31, WPR30, WPR29, WPR28, WPR27, WPR26,
                WPR25, WPR24, WPR23, WPR22, WPR21, WPR20,
                WPR19, WPR18, WPR17, WPR16, WPR15, WPR14,
                WPR13, WPR12, WPR11, WPR10, WPR9,  WPR8,
                WPR7,  WPR6,  WPR5,  WPR4,  WPR3,  WPR2,
                WPR1,  WPR0,*/
		WPR,
		TFCOMPL, RFCOMPL, BUSTMOUT, BUFEND,
		BCNT10, BCNT9,  BCNT8, BCNT7,  BCNT6,  BCNT5,  
		BCNT4,  BCNT3,  BCNT2, BCNT1,  BCNT0,
		TFGNT, RFGNT, BCNTBT40, UMORE, UMORE2LN,
		MBE3_, MBE2_, MBE1_,MBE0_,

		/* input */
		/*BUFPTR31, BUFPTR30, BUFPTR29, BUFPTR28, BUFPTR27, BUFPTR26,
                BUFPTR25, BUFPTR24, BUFPTR23, BUFPTR22, BUFPTR21, BUFPTR20,
                BUFPTR19, BUFPTR18, BUFPTR17, BUFPTR16, BUFPTR15, BUFPTR14,
                BUFPTR13, BUFPTR12, BUFPTR11, BUFPTR10, BUFPTR9,  BUFPTR8,
                BUFPTR7,  BUFPTR6,  BUFPTR5,  BUFPTR4,  BUFPTR3,  BUFPTR2,
                BUFPTR1,  BUFPTR0,*/
		BUFPTR1, BUFPTR2,

		/*MAXLEN10, MAXLEN9,  MAXLEN8, MAXLEN7,  MAXLEN6,  MAXLEN5,  
		MAXLEN4,  MAXLEN3,  MAXLEN2, MAXLEN1,  MAXLEN0,*/
		MAXLEN,
		RFREQ_S, TXREQ, RFLUSH_S,

		FEMPTY, FIFOGNT, PMSTR, RDYACK, 
		/*BUSFREE ,*/NEARFEMP, WPRLD, 
		TXFIFO, RXFIFO, FCFG, 
		/*FBE3_, FBE2_, FBE1_,FBE0_,*/
		FBE_, //UCBE3O_,UCBE2O_,UCBE1O_,UCBE0O_, 
		//PCICLK, PCICLK2, HRST_ 
		PCICLK, HRST_, BOUNDRY, BOUNDRY_T, DIS_BURST, HCIGNT
		);

HS_BMUX HS_BMUX ( 
		/* output */
		//UAD31O, UAD30O, UAD29O, UAD28O, UAD27O, UAD26O,
                //UAD25O, UAD24O, UAD23O, UAD22O, UAD21O, UAD20O,
                //UAD19O, UAD18O, UAD17O, UAD16O, UAD15O, UAD14O,
                //UAD13O, UAD12O, UAD11O, UAD10O, UAD9O,  UAD8O,
                //UAD7O,  UAD6O,  UAD5O,  UAD4O,  UAD3O,  UAD2O,
                //UAD1O,  UAD0O, 

		/* input */
		/*WPR31, WPR30, WPR29, WPR28, WPR27, WPR26,
                WPR25, WPR24, WPR23, WPR22, WPR21, WPR20,
                WPR19, WPR18, WPR17, WPR16, WPR15, WPR14,
                WPR13, WPR12, WPR11, WPR10, WPR9,  WPR8,
                WPR7,  WPR6,  WPR5,  WPR4,  WPR3,  WPR2,
                WPR1,  WPR0,*/
		WPR,

		//PSADO31, PSADO30, PSADO29, PSADO28, PSADO27, PSADO26,
                //PSADO25, PSADO24, PSADO23, PSADO22, PSADO21, PSADO20,
                //PSADO19, PSADO18, PSADO17, PSADO16, PSADO15, PSADO14,
                //PSADO13, PSADO12, PSADO11, PSADO10, PSADO9,  PSADO8,
                //PSADO7,  PSADO6,  PSADO5,  PSADO4,  PSADO3,  PSADO2,
                //PSADO1,  PSADO0,

		/*FFDOUT31, FFDOUT30, FFDOUT29, FFDOUT28, FFDOUT27, FFDOUT26,
                FFDOUT25, FFDOUT24, FFDOUT23, FFDOUT22, FFDOUT21, FFDOUT20,
                FFDOUT19, FFDOUT18, FFDOUT17, FFDOUT16, FFDOUT15, FFDOUT14,
                FFDOUT13, FFDOUT12, FFDOUT11, FFDOUT10, FFDOUT9,  FFDOUT8,
                FFDOUT7,  FFDOUT6,  FFDOUT5,  FFDOUT4,  FFDOUT3,  FFDOUT2,
                FFDOUT1,  FFDOUT0, */
		FFRDPCI,

		/*HCIADR31, HCIADR30, HCIADR29, HCIADR28, HCIADR27, HCIADR26,
                HCIADR25, HCIADR24, HCIADR23, HCIADR22, HCIADR21, HCIADR20,
                HCIADR19, HCIADR18, HCIADR17, HCIADR16, HCIADR15, HCIADR14,
                HCIADR13, HCIADR12, HCIADR11, HCIADR10, HCIADR9,  HCIADR8,
                HCIADR7,  HCIADR6,  HCIADR5,  HCIADR4,  HCIADR3,  HCIADR2,
                HCIADR1,  HCIADR0,
		HCIADD31, HCIADD30, HCIADD29, HCIADD28, HCIADD27, HCIADD26,
                HCIADD25, HCIADD24, HCIADD23, HCIADD22, HCIADD21, HCIADD20,
                HCIADD19, HCIADD18, HCIADD17, HCIADD16, HCIADD15, HCIADD14,
                HCIADD13, HCIADD12, HCIADD11, HCIADD10, HCIADD9,  HCIADD8,
                HCIADD7,  HCIADD6,  HCIADD5,  HCIADD4,  HCIADD3,  HCIADD2,
                HCIADD1,  HCIADD0,*/
		HCIADR, HCIADD,
		/*PMDSEL, PMSTR ,*/ FIFOGNT, HCIGNT,
		MA, MWD
		);

HS_BMUIF HS_BMUIF ( 
		/* output */
		CREQ, MRDY_, CACHEN, COMPL, MSWR, MRDMPLZ, XMITNULL, 
		WPRLD, PCIREAD, PCIWRT, NEARFEMP, NEARFULL, 
		TXTHRESH, RXTHRESH, MYPMACK, //TXTHRESH2, // by Chris Lai

		/* input */
                WPR[1],  WPR[0], BCNTBT40, 
 
		/*MAXLEN10, MAXLEN9,  MAXLEN8, MAXLEN7,  MAXLEN6,  MAXLEN5,  
		MAXLEN4,  MAXLEN3,  MAXLEN2, MAXLEN1,  MAXLEN0,*/
		MAXLEN,

		CACHLN7,  CACHLN6,  CACHLN5,  CACHLN4,  CACHLN3,  CACHLN2,
                CACHLN1,  CACHLN0, CAHCFG_,

		RFCOMPL, TFCOMPL, BUFEND, HCIGNT, FIFOGNT,
		FEMPTY, //FCOUNT4,FCOUNT3,FCOUNT2,FCOUNT1,FCOUNT0, 
		FCOUNT,
		XMITSTRT, RXSTRT, TFGNT, RFGNT, TXREQ, RXREQ,
		/*BUSFREE,*/ RFREQ_S, FCFG, MWRMEN, 
		HCIREQ, HCICOMPL, HCIMWR, HCIMRDY, PMSTR, MADDR, PCI1WAIT, 
		TXFIFO, RXFIFO, EOTQ, RDYACK, PCICLK, HRST_,
		TADOE, /*MADOE,*/ UADOE_, BOUNDRY, BOUNDRY_T, DIS_BURST,
		ZEROLEN, FIFO_OK
		);




// #undef HRST_

endmodule


module HS_DMA_MUX ( MA1, MA2, MA3, MA4, MWD1, MWD2, MWD3, MWD4, MA, MWD, MBE3_, 
    MBE2_, MBE1_, MBE0_, MBE3AI_, MBE2AI_, MBE1AI_, MBE0AI_, MBE3BI_, MBE2BI_, 
    MBE1BI_, MBE0BI_, MBE3CI_, MBE2CI_, MBE1CI_, MBE0CI_, MBE3DI_, MBE2DI_, 
    MBE1DI_, MBE0DI_, CREQ1, CREQ2, CREQ3, CREQ4, CREQ, MRDY1_, MRDY2_, MRDY3_, 
    MRDY4_, MRDY_, CACHEN1, CACHEN2, CACHEN3, CACHEN4, CACHEN, COMPL1, COMPL2, 
    COMPL3, COMPL4, COMPL, MSWR1, MSWR2, MSWR3, MSWR4, MSWR, MRDMPLZ1, 
    MRDMPLZ2, MRDMPLZ3, MRDMPLZ4, MRDMPLZ, HOSTDAT1, HOSTDAT2, HOSTDAT3, 
    HOSTDAT4, HOSTDAT5, HOSTDAT, LATCHDAT1, LATCHDAT2, LATCHDAT3, LATCHDAT4, 
    LATCHDAT5, LATCHDAT, USBPOP1, USBPOP2, USBPOP3, USBPOP4, USBPOP5, USBPOP, 
    BUSFREE1, BUSFREE2, BUSFREE3, BUSFREE4, BUSFREE, UGNTI1_, UGNTI2_, UGNTI3_, 
    UGNTI4_, UGNTI_, PMDSEL1, PMDSEL2, PMDSEL3, PMDSEL4, PMDSEL, PMSTR1, 
    PMSTR2, PMSTR3, PMSTR4, PMSTR, MADDR1, MADDR2, MADDR3, MADDR4, MADDR, 
    RDYACK1, RDYACK2, RDYACK3, RDYACK4, RDYACK, MAXLEN, TRAN_MAXLEN1, 
    SLAVE_ACT, SLAVEMODE, TEST_PACKET, TRAN_BUFPTR1, TRAN_BUFPTR2, DMA_BUFPTR1, 
    DMA_BUFPTR2, SLQUEUEADDR, TXADDR, TXENDP, HUBADDR, HUBPORT, SP_SC, SP_S, 
    SP_E, SP_ET, TD_IN, TD_OUT, TD_SETUP, TD_SPLIT, TD_PING, DAT0, DAT1, DAT2, 
    DATM, ISO, EXEITD, TRAN_CMD1, TRAN_CMD2, TRAN_CMD3, TRAN_CMD4, TRAN_CMD5, 
    PCIDMA_SEL, USBDMA_SEL, BIST_ERR_S1, BIST_ERR_S2, BIST_ERR_S3, BIST_ERR_S4, 
    BIST_ERR_S, UMORE1, UMORE2, UMORE3, UMORE4, UMORE2LN1, UMORE2LN2, 
    UMORE2LN3, UMORE2LN4, UMORE, UMORE2LN, PCICLK, TRST_ );
input  [31:0] MA1;
input  [31:0] MWD2;
input  [31:0] MWD3;
input  [31:0] MWD4;
output [31:0] MA;
input  [7:0] HOSTDAT3;
output [3:0] TXENDP;
output [31:0] DMA_BUFPTR1;
input  [51:0] TRAN_CMD5;
input  [7:0] HOSTDAT4;
output [6:0] HUBPORT;
input  [51:0] TRAN_CMD2;
input  [3:0] PCIDMA_SEL;
output [6:0] TXADDR;
output [31:0] MWD;
input  [7:0] HOSTDAT5;
input  [31:0] TRAN_BUFPTR1;
output [7:0] HOSTDAT;
output [6:0] HUBADDR;
input  [51:0] TRAN_CMD3;
input  [31:0] SLQUEUEADDR;
output [1:0] SP_ET;
input  [4:0] USBDMA_SEL;
input  [31:0] MA2;
input  [31:0] MA3;
input  [7:0] HOSTDAT2;
input  [51:0] TRAN_CMD4;
input  [31:0] MA4;
output [10:0] TRAN_MAXLEN1;
output [19:0] DMA_BUFPTR2;
input  [51:0] TRAN_CMD1;
input  [31:0] MWD1;
input  [19:0] TRAN_BUFPTR2;
output [10:0] MAXLEN;
input  [7:0] HOSTDAT1;
input  MBE3AI_, MBE2AI_, MBE1AI_, MBE0AI_, MBE3BI_, MBE2BI_, MBE1BI_, MBE0BI_, 
    MBE3CI_, MBE2CI_, MBE1CI_, MBE0CI_, MBE3DI_, MBE2DI_, MBE1DI_, MBE0DI_, 
    CREQ1, CREQ2, CREQ3, CREQ4, MRDY1_, MRDY2_, MRDY3_, MRDY4_, CACHEN1, 
    CACHEN2, CACHEN3, CACHEN4, COMPL1, COMPL2, COMPL3, COMPL4, MSWR1, MSWR2, 
    MSWR3, MSWR4, MRDMPLZ1, MRDMPLZ2, MRDMPLZ3, MRDMPLZ4, LATCHDAT, USBPOP, 
    BUSFREE, UGNTI_, PMDSEL, PMSTR, MADDR, RDYACK, SLAVE_ACT, SLAVEMODE, 
    TEST_PACKET, BIST_ERR_S1, BIST_ERR_S2, BIST_ERR_S3, BIST_ERR_S4, UMORE1, 
    UMORE2, UMORE3, UMORE4, UMORE2LN1, UMORE2LN2, UMORE2LN3, UMORE2LN4, PCICLK, 
    TRST_;
output MBE3_, MBE2_, MBE1_, MBE0_, CREQ, MRDY_, CACHEN, COMPL, MSWR, MRDMPLZ, 
    LATCHDAT1, LATCHDAT2, LATCHDAT3, LATCHDAT4, LATCHDAT5, USBPOP1, USBPOP2, 
    USBPOP3, USBPOP4, USBPOP5, BUSFREE1, BUSFREE2, BUSFREE3, BUSFREE4, UGNTI1_, 
    UGNTI2_, UGNTI3_, UGNTI4_, PMDSEL1, PMDSEL2, PMDSEL3, PMDSEL4, PMSTR1, 
    PMSTR2, PMSTR3, PMSTR4, MADDR1, MADDR2, MADDR3, MADDR4, RDYACK1, RDYACK2, 
    RDYACK3, RDYACK4, SP_SC, SP_S, SP_E, TD_IN, TD_OUT, TD_SETUP, TD_SPLIT, 
    TD_PING, DAT0, DAT1, DAT2, DATM, ISO, EXEITD, BIST_ERR_S, UMORE, UMORE2LN;
    wire b997_19, SPAREO6, b997_9, b997_10, SPAREO0_, b997_7, b997_17, SPAREO8, 
        SPAREO1, b997_16, SPAREO9, b997_6, SPAREO0, b997_8, b997_18, SPAREO7, 
        b997_11, SPAREO5, b997_13, b997_3, b997_4, b997_14, SPAREO2, b997_15, 
        b997_5, SPAREO3, SPAREO1_, SPAREO4, b997_2, b997_12, n1148, n1149, 
        n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
        n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
        n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
        n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
        n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
        n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
        n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
        n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
        n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
        n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
        n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
        n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
        n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
        n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
        n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
        n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
        n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
        n1320, n1321, n1322, n1323, n1324, n1325, n1326, add_231_carry_15, 
        add_231_carry_8, add_231_carry_12, add_231_carry_6, add_231_carry_14, 
        add_231_carry_13, add_231_carry_7, add_231_carry_16, add_231_carry_9, 
        add_231_carry_2, add_231_carry_18, add_231_carry_11, add_231_carry_5, 
        add_231_carry_19, add_231_carry_4, add_231_carry_10, add_231_carry_17, 
        add_231_carry_3;
    zaoi211b SPARE822 ( .A(SPAREO0), .B(1'b1), .C(SPAREO1_), .D(1'b0), .Y(
        SPAREO2) );
    zoai21b SPARE825 ( .A(SPAREO1), .B(1'b0), .C(SPAREO9), .Y(SPAREO3) );
    zoai21b SPARE824 ( .A(SPAREO0), .B(SPAREO8), .C(1'b1), .Y(SPAREO9) );
    zaoi211b SPARE823 ( .A(SPAREO4), .B(1'b1), .C(SPAREO6), .D(1'b0), .Y(
        SPAREO8) );
    zdffrb SPARE821 ( .CK(PCICLK), .D(SPAREO7), .R(TRST_), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE828 ( .A(SPAREO5), .Y(SPAREO6) );
    znr3b SPARE826 ( .A(SPAREO2), .B(MSWR), .C(SPAREO0_), .Y(SPAREO4) );
    zivb SPARE827 ( .A(SPAREO4), .Y(SPAREO5) );
    zdffrb SPARE820 ( .CK(PCICLK), .D(1'b0), .R(TRST_), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE829 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zhadrb add_231_U1_1_1 ( .A(SLQUEUEADDR[13]), .B(SLQUEUEADDR[12]), .CO(
        add_231_carry_2), .S(b997_2) );
    zhadrb add_231_U1_1_2 ( .A(SLQUEUEADDR[14]), .B(add_231_carry_2), .CO(
        add_231_carry_3), .S(b997_3) );
    zhadrb add_231_U1_1_3 ( .A(SLQUEUEADDR[15]), .B(add_231_carry_3), .CO(
        add_231_carry_4), .S(b997_4) );
    zhadrb add_231_U1_1_4 ( .A(SLQUEUEADDR[16]), .B(add_231_carry_4), .CO(
        add_231_carry_5), .S(b997_5) );
    zhadrb add_231_U1_1_5 ( .A(SLQUEUEADDR[17]), .B(add_231_carry_5), .CO(
        add_231_carry_6), .S(b997_6) );
    zhadrb add_231_U1_1_6 ( .A(SLQUEUEADDR[18]), .B(add_231_carry_6), .CO(
        add_231_carry_7), .S(b997_7) );
    zhadrb add_231_U1_1_7 ( .A(SLQUEUEADDR[19]), .B(add_231_carry_7), .CO(
        add_231_carry_8), .S(b997_8) );
    zhadrb add_231_U1_1_8 ( .A(SLQUEUEADDR[20]), .B(add_231_carry_8), .CO(
        add_231_carry_9), .S(b997_9) );
    zhadrb add_231_U1_1_9 ( .A(SLQUEUEADDR[21]), .B(add_231_carry_9), .CO(
        add_231_carry_10), .S(b997_10) );
    zhadrb add_231_U1_1_10 ( .A(SLQUEUEADDR[22]), .B(add_231_carry_10), .CO(
        add_231_carry_11), .S(b997_11) );
    zhadrb add_231_U1_1_11 ( .A(SLQUEUEADDR[23]), .B(add_231_carry_11), .CO(
        add_231_carry_12), .S(b997_12) );
    zhadrb add_231_U1_1_12 ( .A(SLQUEUEADDR[24]), .B(add_231_carry_12), .CO(
        add_231_carry_13), .S(b997_13) );
    zhadrb add_231_U1_1_13 ( .A(SLQUEUEADDR[25]), .B(add_231_carry_13), .CO(
        add_231_carry_14), .S(b997_14) );
    zhadrb add_231_U1_1_14 ( .A(SLQUEUEADDR[26]), .B(add_231_carry_14), .CO(
        add_231_carry_15), .S(b997_15) );
    zhadrb add_231_U1_1_15 ( .A(SLQUEUEADDR[27]), .B(add_231_carry_15), .CO(
        add_231_carry_16), .S(b997_16) );
    zhadrb add_231_U1_1_16 ( .A(SLQUEUEADDR[28]), .B(add_231_carry_16), .CO(
        add_231_carry_17), .S(b997_17) );
    zhadrb add_231_U1_1_17 ( .A(SLQUEUEADDR[29]), .B(add_231_carry_17), .CO(
        add_231_carry_18), .S(b997_18) );
    zhadrb add_231_U1_1_18 ( .A(SLQUEUEADDR[30]), .B(add_231_carry_18), .CO(
        add_231_carry_19), .S(b997_19) );
    zivb U90 ( .A(n1185), .Y(n1148) );
    zivb U91 ( .A(n1178), .Y(n1150) );
    zivb U92 ( .A(n1178), .Y(n1149) );
    zivb U93 ( .A(n1178), .Y(n1195) );
    zbfb U94 ( .A(n1323), .Y(n1151) );
    zbfb U95 ( .A(n1323), .Y(n1153) );
    zbfb U96 ( .A(n1323), .Y(n1152) );
    znd3b U97 ( .A(n1320), .B(n1180), .C(USBDMA_SEL[2]), .Y(n1154) );
    zivb U98 ( .A(n1154), .Y(n1155) );
    zivb U99 ( .A(n1154), .Y(n1157) );
    zivb U100 ( .A(n1154), .Y(n1156) );
    zivb U101 ( .A(n1213), .Y(n1158) );
    zivb U102 ( .A(n1158), .Y(n1159) );
    zivb U103 ( .A(n1158), .Y(n1162) );
    zivb U104 ( .A(n1158), .Y(n1160) );
    zivb U105 ( .A(n1158), .Y(n1161) );
    zivb U106 ( .A(n1214), .Y(n1163) );
    zivb U107 ( .A(n1163), .Y(n1164) );
    zivb U108 ( .A(n1163), .Y(n1167) );
    zivb U109 ( .A(n1163), .Y(n1165) );
    zivb U110 ( .A(n1163), .Y(n1166) );
    znd2b U111 ( .A(PCIDMA_SEL[2]), .B(n1321), .Y(n1168) );
    zivb U112 ( .A(n1168), .Y(n1169) );
    zivb U113 ( .A(n1168), .Y(n1172) );
    zivb U114 ( .A(n1168), .Y(n1170) );
    zivb U115 ( .A(n1168), .Y(n1171) );
    zor2b U116 ( .A(USBDMA_SEL[3]), .B(n1322), .Y(n1173) );
    zivb U117 ( .A(n1173), .Y(n1174) );
    zivb U118 ( .A(n1173), .Y(n1176) );
    zivb U119 ( .A(n1173), .Y(n1175) );
    zbfb U120 ( .A(SLAVEMODE), .Y(n1177) );
    zbfb U121 ( .A(SLAVEMODE), .Y(n1179) );
    zbfb U122 ( .A(SLAVEMODE), .Y(n1178) );
    zivb U123 ( .A(USBDMA_SEL[0]), .Y(n1180) );
    zivb U124 ( .A(n1180), .Y(n1181) );
    zivb U125 ( .A(n1180), .Y(n1184) );
    zivb U126 ( .A(n1180), .Y(n1182) );
    zivb U127 ( .A(n1180), .Y(n1183) );
    zivb U128 ( .A(PCIDMA_SEL[0]), .Y(n1185) );
    zivb U129 ( .A(n1185), .Y(n1186) );
    zivb U130 ( .A(n1185), .Y(n1189) );
    zivb U131 ( .A(n1185), .Y(n1187) );
    zivb U132 ( .A(n1185), .Y(n1188) );
    zinr2d U133 ( .A(USBDMA_SEL[3]), .B(n1322), .Y(n1323) );
    zinr2d U134 ( .A(n1321), .B(PCIDMA_SEL[2]), .Y(n1213) );
    zinr2d U135 ( .A(PCIDMA_SEL[1]), .B(n1189), .Y(n1214) );
    zor2b U136 ( .A(n1183), .B(n1320), .Y(n1190) );
    zivb U137 ( .A(n1190), .Y(n1191) );
    zivb U138 ( .A(n1190), .Y(n1193) );
    zivb U139 ( .A(n1190), .Y(n1192) );
    zao21b U140 ( .A(TRAN_CMD1[50]), .B(n1194), .C(n1178), .Y(TRAN_MAXLEN1[10]
        ) );
    zao21b U141 ( .A(TRAN_CMD1[45]), .B(n1195), .C(n1196), .Y(TRAN_MAXLEN1[5])
         );
    zao21b U142 ( .A(TRAN_CMD1[44]), .B(n1195), .C(n1196), .Y(TRAN_MAXLEN1[4])
         );
    zao21b U143 ( .A(TRAN_CMD1[42]), .B(n1150), .C(n1196), .Y(TRAN_MAXLEN1[2])
         );
    zao21b U144 ( .A(TRAN_CMD1[40]), .B(n1150), .C(n1196), .Y(TRAN_MAXLEN1[0])
         );
    zao21b U145 ( .A(n1197), .B(n1194), .C(n1178), .Y(MAXLEN[10]) );
    zao22b U146 ( .A(TRAN_MAXLEN1[9]), .B(n1181), .C(n1198), .D(n1199), .Y(
        MAXLEN[9]) );
    zao22b U147 ( .A(TRAN_MAXLEN1[8]), .B(n1184), .C(n1198), .D(n1200), .Y(
        MAXLEN[8]) );
    zao22b U148 ( .A(TRAN_MAXLEN1[7]), .B(n1183), .C(n1198), .D(n1201), .Y(
        MAXLEN[7]) );
    zao22b U149 ( .A(TRAN_MAXLEN1[6]), .B(n1184), .C(n1198), .D(n1202), .Y(
        MAXLEN[6]) );
    zoa21b U150 ( .A(n1203), .B(n1204), .C(n1195), .Y(MAXLEN[5]) );
    zoa21b U151 ( .A(n1205), .B(n1206), .C(n1150), .Y(MAXLEN[4]) );
    zao22b U152 ( .A(TRAN_MAXLEN1[3]), .B(n1182), .C(n1198), .D(n1207), .Y(
        MAXLEN[3]) );
    zoa21b U153 ( .A(n1208), .B(n1209), .C(n1195), .Y(MAXLEN[2]) );
    zao22b U154 ( .A(TRAN_MAXLEN1[1]), .B(n1181), .C(n1198), .D(n1210), .Y(
        MAXLEN[1]) );
    zoa21b U155 ( .A(n1211), .B(n1212), .C(n1150), .Y(MAXLEN[0]) );
    zao2x4b U156 ( .A(MA1[0]), .B(n1188), .C(MA3[0]), .D(n1170), .E(MA4[0]), 
        .F(n1160), .G(MA2[0]), .H(n1166), .Y(MA[0]) );
    zao2x4b U157 ( .A(MA1[1]), .B(n1187), .C(MA3[1]), .D(n1170), .E(MA4[1]), 
        .F(n1162), .G(MA2[1]), .H(n1164), .Y(MA[1]) );
    zao2x4b U158 ( .A(MA1[2]), .B(n1189), .C(MA3[2]), .D(n1170), .E(MA4[2]), 
        .F(n1160), .G(MA2[2]), .H(n1166), .Y(MA[2]) );
    zao2x4b U159 ( .A(MA1[3]), .B(n1148), .C(MA3[3]), .D(n1169), .E(MA4[3]), 
        .F(n1159), .G(MA2[3]), .H(n1164), .Y(MA[3]) );
    zao2x4b U160 ( .A(MA1[4]), .B(n1189), .C(MA3[4]), .D(n1171), .E(MA4[4]), 
        .F(n1161), .G(MA2[4]), .H(n1166), .Y(MA[4]) );
    zao2x4b U161 ( .A(MA1[5]), .B(n1187), .C(MA3[5]), .D(n1171), .E(MA4[5]), 
        .F(n1162), .G(MA2[5]), .H(n1164), .Y(MA[5]) );
    zao2x4b U162 ( .A(MA1[6]), .B(n1187), .C(MA3[6]), .D(n1172), .E(MA4[6]), 
        .F(n1160), .G(MA2[6]), .H(n1166), .Y(MA[6]) );
    zao2x4b U163 ( .A(MA1[7]), .B(n1189), .C(MA3[7]), .D(n1169), .E(MA4[7]), 
        .F(n1162), .G(MA2[7]), .H(n1167), .Y(MA[7]) );
    zao2x4b U164 ( .A(MA1[8]), .B(n1187), .C(MA3[8]), .D(n1171), .E(MA4[8]), 
        .F(n1160), .G(MA2[8]), .H(n1165), .Y(MA[8]) );
    zao2x4b U165 ( .A(MA1[9]), .B(n1186), .C(MA3[9]), .D(n1170), .E(MA4[9]), 
        .F(n1159), .G(MA2[9]), .H(n1164), .Y(MA[9]) );
    zao2x4b U166 ( .A(MA1[10]), .B(n1188), .C(MA3[10]), .D(n1170), .E(MA4[10]), 
        .F(n1161), .G(MA2[10]), .H(n1166), .Y(MA[10]) );
    zao2x4b U167 ( .A(MA1[11]), .B(n1188), .C(MA3[11]), .D(n1170), .E(MA4[11]), 
        .F(n1159), .G(MA2[11]), .H(n1164), .Y(MA[11]) );
    zao2x4b U168 ( .A(MA1[12]), .B(n1187), .C(MA3[12]), .D(n1171), .E(MA4[12]), 
        .F(n1161), .G(MA2[12]), .H(n1166), .Y(MA[12]) );
    zao2x4b U169 ( .A(MA1[13]), .B(n1186), .C(MA3[13]), .D(n1171), .E(MA4[13]), 
        .F(n1159), .G(MA2[13]), .H(n1164), .Y(MA[13]) );
    zao2x4b U170 ( .A(MA1[14]), .B(n1148), .C(MA3[14]), .D(n1172), .E(MA4[14]), 
        .F(n1161), .G(MA2[14]), .H(n1166), .Y(MA[14]) );
    zao2x4b U171 ( .A(MA1[15]), .B(n1148), .C(MA3[15]), .D(n1170), .E(MA4[15]), 
        .F(n1162), .G(MA2[15]), .H(n1164), .Y(MA[15]) );
    zao2x4b U172 ( .A(MA1[16]), .B(n1188), .C(MA3[16]), .D(n1171), .E(MA4[16]), 
        .F(n1160), .G(MA2[16]), .H(n1166), .Y(MA[16]) );
    zao2x4b U173 ( .A(MA1[17]), .B(n1188), .C(MA3[17]), .D(n1171), .E(MA4[17]), 
        .F(n1162), .G(MA2[17]), .H(n1167), .Y(MA[17]) );
    zao2x4b U174 ( .A(MA1[18]), .B(n1186), .C(MA3[18]), .D(n1172), .E(MA4[18]), 
        .F(n1160), .G(MA2[18]), .H(n1165), .Y(MA[18]) );
    zao2x4b U175 ( .A(MA1[19]), .B(n1186), .C(MA3[19]), .D(n1170), .E(MA4[19]), 
        .F(n1162), .G(MA2[19]), .H(n1167), .Y(MA[19]) );
    zao2x4b U176 ( .A(MA1[20]), .B(n1186), .C(MA3[20]), .D(n1171), .E(MA4[20]), 
        .F(n1160), .G(MA2[20]), .H(n1165), .Y(MA[20]) );
    zao2x4b U177 ( .A(MA1[21]), .B(n1188), .C(MA3[21]), .D(n1170), .E(MA4[21]), 
        .F(n1162), .G(MA2[21]), .H(n1167), .Y(MA[21]) );
    zao2x4b U178 ( .A(MA1[22]), .B(n1187), .C(MA3[22]), .D(n1172), .E(MA4[22]), 
        .F(n1160), .G(MA2[22]), .H(n1165), .Y(MA[22]) );
    zao2x4b U179 ( .A(MA1[23]), .B(n1187), .C(MA3[23]), .D(n1170), .E(MA4[23]), 
        .F(n1162), .G(MA2[23]), .H(n1167), .Y(MA[23]) );
    zao2x4b U180 ( .A(MA1[24]), .B(n1189), .C(MA3[24]), .D(n1170), .E(MA4[24]), 
        .F(n1160), .G(MA2[24]), .H(n1165), .Y(MA[24]) );
    zao2x4b U181 ( .A(MA1[25]), .B(n1189), .C(MA3[25]), .D(n1171), .E(MA4[25]), 
        .F(n1162), .G(MA2[25]), .H(n1167), .Y(MA[25]) );
    zao2x4b U182 ( .A(MA1[26]), .B(n1189), .C(MA3[26]), .D(n1171), .E(MA4[26]), 
        .F(n1160), .G(MA2[26]), .H(n1165), .Y(MA[26]) );
    zao2x4b U183 ( .A(MA1[27]), .B(n1148), .C(MA3[27]), .D(n1169), .E(MA4[27]), 
        .F(n1162), .G(MA2[27]), .H(n1164), .Y(MA[27]) );
    zao2x4b U184 ( .A(MA1[28]), .B(n1148), .C(MA3[28]), .D(n1171), .E(MA4[28]), 
        .F(n1160), .G(MA2[28]), .H(n1166), .Y(MA[28]) );
    zao2x4b U185 ( .A(MA1[29]), .B(n1186), .C(MA3[29]), .D(n1170), .E(MA4[29]), 
        .F(n1162), .G(MA2[29]), .H(n1167), .Y(MA[29]) );
    zao2x4b U186 ( .A(MA1[30]), .B(n1189), .C(MA3[30]), .D(n1172), .E(MA4[30]), 
        .F(n1160), .G(MA2[30]), .H(n1165), .Y(MA[30]) );
    zao2x4b U187 ( .A(MA1[31]), .B(n1187), .C(MA3[31]), .D(n1171), .E(MA4[31]), 
        .F(n1162), .G(MA2[31]), .H(n1167), .Y(MA[31]) );
    zao2x4b U188 ( .A(MBE0AI_), .B(n1188), .C(MBE0CI_), .D(n1171), .E(MBE0DI_), 
        .F(n1160), .G(MBE0BI_), .H(n1165), .Y(MBE0_) );
    zao2x4b U189 ( .A(MBE1AI_), .B(n1148), .C(MBE1CI_), .D(n1171), .E(MBE1DI_), 
        .F(n1162), .G(MBE1BI_), .H(n1167), .Y(MBE1_) );
    zao2x4b U190 ( .A(MBE2AI_), .B(n1187), .C(MBE2CI_), .D(n1171), .E(MBE2DI_), 
        .F(n1160), .G(MBE2BI_), .H(n1165), .Y(MBE2_) );
    zao2x4b U191 ( .A(MBE3AI_), .B(n1148), .C(MBE3CI_), .D(n1170), .E(MBE3DI_), 
        .F(n1159), .G(MBE3BI_), .H(n1164), .Y(MBE3_) );
    zao211b U192 ( .A(TRAN_CMD3[1]), .B(n1157), .C(n1215), .D(n1216), .Y(DATM)
         );
    zao211b U193 ( .A(TRAN_CMD3[2]), .B(n1156), .C(n1217), .D(n1218), .Y(DAT2)
         );
    zao211b U194 ( .A(TRAN_CMD3[3]), .B(n1156), .C(n1219), .D(n1220), .Y(DAT1)
         );
    zao211b U195 ( .A(TRAN_CMD3[4]), .B(n1156), .C(n1221), .D(n1222), .Y(DAT0)
         );
    zao211b U196 ( .A(TRAN_CMD3[5]), .B(n1155), .C(n1223), .D(n1224), .Y(
        TD_PING) );
    zao211b U197 ( .A(TRAN_CMD3[6]), .B(n1155), .C(n1225), .D(n1226), .Y(
        TD_SPLIT) );
    zao211b U198 ( .A(TRAN_CMD3[7]), .B(n1155), .C(n1227), .D(n1228), .Y(
        TD_SETUP) );
    zao211b U199 ( .A(TRAN_CMD3[8]), .B(n1156), .C(n1229), .D(n1230), .Y(
        TD_OUT) );
    zao211b U200 ( .A(TRAN_CMD3[9]), .B(n1155), .C(n1231), .D(n1232), .Y(TD_IN
        ) );
    zao211b U201 ( .A(TRAN_CMD3[10]), .B(n1157), .C(n1233), .D(n1234), .Y(
        SP_ET[0]) );
    zao211b U202 ( .A(TRAN_CMD3[11]), .B(n1157), .C(n1235), .D(n1236), .Y(
        SP_ET[1]) );
    zao211b U203 ( .A(TRAN_CMD3[12]), .B(n1157), .C(n1237), .D(n1238), .Y(SP_E
        ) );
    zao211b U204 ( .A(TRAN_CMD3[13]), .B(n1156), .C(n1239), .D(n1240), .Y(SP_S
        ) );
    zao211b U205 ( .A(TRAN_CMD3[14]), .B(n1156), .C(n1241), .D(n1242), .Y(
        SP_SC) );
    zao211b U206 ( .A(TRAN_CMD3[15]), .B(n1155), .C(n1243), .D(n1244), .Y(
        HUBPORT[0]) );
    zao211b U207 ( .A(TRAN_CMD3[16]), .B(n1155), .C(n1245), .D(n1246), .Y(
        HUBPORT[1]) );
    zao211b U208 ( .A(TRAN_CMD3[17]), .B(n1156), .C(n1247), .D(n1248), .Y(
        HUBPORT[2]) );
    zao211b U209 ( .A(TRAN_CMD3[18]), .B(n1155), .C(n1249), .D(n1250), .Y(
        HUBPORT[3]) );
    zao211b U210 ( .A(TRAN_CMD3[19]), .B(n1156), .C(n1251), .D(n1252), .Y(
        HUBPORT[4]) );
    zao211b U211 ( .A(TRAN_CMD3[20]), .B(n1156), .C(n1253), .D(n1254), .Y(
        HUBPORT[5]) );
    zao211b U212 ( .A(TRAN_CMD3[21]), .B(n1157), .C(n1255), .D(n1256), .Y(
        HUBPORT[6]) );
    zao211b U213 ( .A(TRAN_CMD3[22]), .B(n1157), .C(n1257), .D(n1258), .Y(
        HUBADDR[0]) );
    zao211b U214 ( .A(TRAN_CMD3[23]), .B(n1157), .C(n1259), .D(n1260), .Y(
        HUBADDR[1]) );
    zao211b U215 ( .A(TRAN_CMD3[24]), .B(n1156), .C(n1261), .D(n1262), .Y(
        HUBADDR[2]) );
    zao211b U216 ( .A(TRAN_CMD3[25]), .B(n1157), .C(n1263), .D(n1264), .Y(
        HUBADDR[3]) );
    zao211b U217 ( .A(TRAN_CMD3[26]), .B(n1157), .C(n1265), .D(n1266), .Y(
        HUBADDR[4]) );
    zao211b U218 ( .A(TRAN_CMD3[27]), .B(n1155), .C(n1267), .D(n1268), .Y(
        HUBADDR[5]) );
    zao211b U219 ( .A(TRAN_CMD3[28]), .B(n1156), .C(n1269), .D(n1270), .Y(
        HUBADDR[6]) );
    zao211b U220 ( .A(TRAN_CMD3[29]), .B(n1156), .C(n1271), .D(n1272), .Y(
        TXENDP[0]) );
    zao211b U221 ( .A(TRAN_CMD3[30]), .B(n1155), .C(n1273), .D(n1274), .Y(
        TXENDP[1]) );
    zao211b U222 ( .A(TRAN_CMD3[31]), .B(n1157), .C(n1275), .D(n1276), .Y(
        TXENDP[2]) );
    zao211b U223 ( .A(TRAN_CMD3[32]), .B(n1155), .C(n1277), .D(n1278), .Y(
        TXENDP[3]) );
    zao211b U224 ( .A(TRAN_CMD3[33]), .B(n1157), .C(n1279), .D(n1280), .Y(
        TXADDR[0]) );
    zao211b U225 ( .A(TRAN_CMD3[34]), .B(n1155), .C(n1281), .D(n1282), .Y(
        TXADDR[1]) );
    zao211b U226 ( .A(TRAN_CMD3[35]), .B(n1157), .C(n1283), .D(n1284), .Y(
        TXADDR[2]) );
    zao211b U227 ( .A(TRAN_CMD3[36]), .B(n1156), .C(n1285), .D(n1286), .Y(
        TXADDR[3]) );
    zao211b U228 ( .A(TRAN_CMD3[37]), .B(n1155), .C(n1287), .D(n1288), .Y(
        TXADDR[4]) );
    zao211b U229 ( .A(TRAN_CMD3[38]), .B(n1156), .C(n1289), .D(n1290), .Y(
        TXADDR[5]) );
    zao211b U230 ( .A(TRAN_CMD3[39]), .B(n1157), .C(n1291), .D(n1292), .Y(
        TXADDR[6]) );
    zao211b U231 ( .A(TRAN_CMD3[51]), .B(n1155), .C(n1293), .D(n1294), .Y(
        EXEITD) );
    zao2x4b U232 ( .A(MWD1[0]), .B(n1186), .C(MWD3[0]), .D(n1171), .E(MWD4[0]), 
        .F(n1161), .G(MWD2[0]), .H(n1166), .Y(MWD[0]) );
    zao2x4b U233 ( .A(MWD1[1]), .B(n1189), .C(MWD3[1]), .D(n1169), .E(MWD4[1]), 
        .F(n1160), .G(MWD2[1]), .H(n1165), .Y(MWD[1]) );
    zao2x4b U234 ( .A(MWD1[2]), .B(n1148), .C(MWD3[2]), .D(n1170), .E(MWD4[2]), 
        .F(n1159), .G(MWD2[2]), .H(n1164), .Y(MWD[2]) );
    zao2x4b U235 ( .A(MWD1[3]), .B(n1189), .C(MWD3[3]), .D(n1172), .E(MWD4[3]), 
        .F(n1162), .G(MWD2[3]), .H(n1167), .Y(MWD[3]) );
    zao2x4b U236 ( .A(MWD1[4]), .B(n1188), .C(MWD3[4]), .D(n1172), .E(MWD4[4]), 
        .F(n1161), .G(MWD2[4]), .H(n1166), .Y(MWD[4]) );
    zao2x4b U237 ( .A(MWD1[5]), .B(n1187), .C(MWD3[5]), .D(n1172), .E(MWD4[5]), 
        .F(n1159), .G(MWD2[5]), .H(n1165), .Y(MWD[5]) );
    zao2x4b U238 ( .A(MWD1[6]), .B(n1186), .C(MWD3[6]), .D(n1169), .E(MWD4[6]), 
        .F(n1159), .G(MWD2[6]), .H(n1164), .Y(MWD[6]) );
    zao2x4b U239 ( .A(MWD1[7]), .B(n1148), .C(MWD3[7]), .D(n1170), .E(MWD4[7]), 
        .F(n1160), .G(MWD2[7]), .H(n1165), .Y(MWD[7]) );
    zao2x4b U240 ( .A(MWD1[8]), .B(n1186), .C(MWD3[8]), .D(n1172), .E(MWD4[8]), 
        .F(n1161), .G(MWD2[8]), .H(n1166), .Y(MWD[8]) );
    zao2x4b U241 ( .A(MWD1[9]), .B(n1187), .C(MWD3[9]), .D(n1172), .E(MWD4[9]), 
        .F(n1161), .G(MWD2[9]), .H(n1167), .Y(MWD[9]) );
    zao2x4b U242 ( .A(MWD1[10]), .B(n1148), .C(MWD3[10]), .D(n1171), .E(MWD4
        [10]), .F(n1159), .G(MWD2[10]), .H(n1164), .Y(MWD[10]) );
    zao2x4b U243 ( .A(MWD1[11]), .B(n1148), .C(MWD3[11]), .D(n1170), .E(MWD4
        [11]), .F(n1162), .G(MWD2[11]), .H(n1167), .Y(MWD[11]) );
    zao2x4b U244 ( .A(MWD1[12]), .B(n1188), .C(MWD3[12]), .D(n1170), .E(MWD4
        [12]), .F(n1161), .G(MWD2[12]), .H(n1166), .Y(MWD[12]) );
    zao2x4b U245 ( .A(MWD1[13]), .B(n1148), .C(MWD3[13]), .D(n1172), .E(MWD4
        [13]), .F(n1161), .G(MWD2[13]), .H(n1167), .Y(MWD[13]) );
    zao2x4b U246 ( .A(MWD1[14]), .B(n1189), .C(MWD3[14]), .D(n1169), .E(MWD4
        [14]), .F(n1159), .G(MWD2[14]), .H(n1164), .Y(MWD[14]) );
    zao2x4b U247 ( .A(MWD1[15]), .B(n1186), .C(MWD3[15]), .D(n1171), .E(MWD4
        [15]), .F(n1160), .G(MWD2[15]), .H(n1165), .Y(MWD[15]) );
    zao2x4b U248 ( .A(MWD1[16]), .B(n1187), .C(MWD3[16]), .D(n1172), .E(MWD4
        [16]), .F(n1161), .G(MWD2[16]), .H(n1166), .Y(MWD[16]) );
    zao2x4b U249 ( .A(MWD1[17]), .B(n1188), .C(MWD3[17]), .D(n1172), .E(MWD4
        [17]), .F(n1159), .G(MWD2[17]), .H(n1165), .Y(MWD[17]) );
    zao2x4b U250 ( .A(MWD1[18]), .B(n1186), .C(MWD3[18]), .D(n1169), .E(MWD4
        [18]), .F(n1159), .G(MWD2[18]), .H(n1164), .Y(MWD[18]) );
    zao2x4b U251 ( .A(MWD1[19]), .B(n1188), .C(MWD3[19]), .D(n1172), .E(MWD4
        [19]), .F(n1162), .G(MWD2[19]), .H(n1167), .Y(MWD[19]) );
    zao2x4b U252 ( .A(MWD1[20]), .B(n1189), .C(MWD3[20]), .D(n1169), .E(MWD4
        [20]), .F(n1161), .G(MWD2[20]), .H(n1167), .Y(MWD[20]) );
    zao2x4b U253 ( .A(MWD1[21]), .B(n1188), .C(MWD3[21]), .D(n1169), .E(MWD4
        [21]), .F(n1162), .G(MWD2[21]), .H(n1167), .Y(MWD[21]) );
    zao2x4b U254 ( .A(MWD1[22]), .B(n1148), .C(MWD3[22]), .D(n1169), .E(MWD4
        [22]), .F(n1159), .G(MWD2[22]), .H(n1165), .Y(MWD[22]) );
    zao2x4b U255 ( .A(MWD1[23]), .B(n1187), .C(MWD3[23]), .D(n1169), .E(MWD4
        [23]), .F(n1160), .G(MWD2[23]), .H(n1165), .Y(MWD[23]) );
    zao2x4b U256 ( .A(MWD1[24]), .B(n1148), .C(MWD3[24]), .D(n1169), .E(MWD4
        [24]), .F(n1161), .G(MWD2[24]), .H(n1166), .Y(MWD[24]) );
    zao2x4b U257 ( .A(MWD1[25]), .B(n1186), .C(MWD3[25]), .D(n1169), .E(MWD4
        [25]), .F(n1161), .G(MWD2[25]), .H(n1166), .Y(MWD[25]) );
    zao2x4b U258 ( .A(MWD1[26]), .B(n1186), .C(MWD3[26]), .D(n1172), .E(MWD4
        [26]), .F(n1159), .G(MWD2[26]), .H(n1164), .Y(MWD[26]) );
    zao2x4b U259 ( .A(MWD1[27]), .B(n1188), .C(MWD3[27]), .D(n1169), .E(MWD4
        [27]), .F(n1161), .G(MWD2[27]), .H(n1167), .Y(MWD[27]) );
    zao2x4b U260 ( .A(MWD1[28]), .B(n1189), .C(MWD3[28]), .D(n1172), .E(MWD4
        [28]), .F(n1161), .G(MWD2[28]), .H(n1166), .Y(MWD[28]) );
    zao2x4b U261 ( .A(MWD1[29]), .B(n1186), .C(MWD3[29]), .D(n1169), .E(MWD4
        [29]), .F(n1159), .G(MWD2[29]), .H(n1165), .Y(MWD[29]) );
    zao2x4b U262 ( .A(MWD1[30]), .B(n1148), .C(MWD3[30]), .D(n1169), .E(MWD4
        [30]), .F(n1159), .G(MWD2[30]), .H(n1164), .Y(MWD[30]) );
    zao2x4b U263 ( .A(MWD1[31]), .B(n1189), .C(MWD3[31]), .D(n1172), .E(MWD4
        [31]), .F(n1159), .G(MWD2[31]), .H(n1165), .Y(MWD[31]) );
    zao211b U264 ( .A(HOSTDAT3[0]), .B(n1156), .C(n1295), .D(n1296), .Y(
        HOSTDAT[0]) );
    zao211b U265 ( .A(HOSTDAT3[1]), .B(n1157), .C(n1297), .D(n1298), .Y(
        HOSTDAT[1]) );
    zao211b U266 ( .A(HOSTDAT3[2]), .B(n1157), .C(n1299), .D(n1300), .Y(
        HOSTDAT[2]) );
    zao211b U267 ( .A(HOSTDAT3[3]), .B(n1155), .C(n1301), .D(n1302), .Y(
        HOSTDAT[3]) );
    zao211b U268 ( .A(HOSTDAT3[4]), .B(n1156), .C(n1303), .D(n1304), .Y(
        HOSTDAT[4]) );
    zao211b U269 ( .A(HOSTDAT3[5]), .B(n1155), .C(n1305), .D(n1306), .Y(
        HOSTDAT[5]) );
    zao211b U270 ( .A(HOSTDAT3[6]), .B(n1155), .C(n1307), .D(n1308), .Y(
        HOSTDAT[6]) );
    zao211b U271 ( .A(HOSTDAT3[7]), .B(n1156), .C(n1309), .D(n1310), .Y(
        HOSTDAT[7]) );
    zao2x4b U272 ( .A(UMORE1), .B(n1188), .C(UMORE3), .D(n1170), .E(UMORE4), 
        .F(n1161), .G(UMORE2), .H(n1166), .Y(UMORE) );
    zao2x4b U273 ( .A(n1187), .B(UMORE2LN1), .C(UMORE2LN3), .D(n1169), .E(
        UMORE2LN4), .F(n1159), .G(UMORE2LN2), .H(n1164), .Y(UMORE2LN) );
    zan2b U274 ( .A(MADDR), .B(PCIDMA_SEL[2]), .Y(MADDR3) );
    zan2b U275 ( .A(LATCHDAT), .B(USBDMA_SEL[2]), .Y(LATCHDAT3) );
    zoa21b U276 ( .A(n1311), .B(n1312), .C(n1313), .Y(ISO) );
    znd2b U277 ( .A(PCIDMA_SEL[2]), .B(n1314), .Y(UGNTI3_) );
    znd2b U278 ( .A(PCIDMA_SEL[3]), .B(n1314), .Y(UGNTI4_) );
    zan2b U279 ( .A(USBPOP), .B(USBDMA_SEL[4]), .Y(USBPOP5) );
    zan2b U280 ( .A(MADDR), .B(n1187), .Y(MADDR1) );
    zao2x4b U281 ( .A(CACHEN1), .B(n1189), .C(CACHEN3), .D(PCIDMA_SEL[2]), .E(
        CACHEN4), .F(PCIDMA_SEL[3]), .G(CACHEN2), .H(PCIDMA_SEL[1]), .Y(CACHEN
        ) );
    zan2b U282 ( .A(PMSTR), .B(PCIDMA_SEL[3]), .Y(PMSTR4) );
    zan2b U283 ( .A(BUSFREE), .B(PCIDMA_SEL[1]), .Y(BUSFREE2) );
    zan2b U284 ( .A(RDYACK), .B(PCIDMA_SEL[3]), .Y(RDYACK4) );
    zan2b U285 ( .A(USBDMA_SEL[3]), .B(USBPOP), .Y(USBPOP4) );
    zan2b U286 ( .A(PMDSEL), .B(n1186), .Y(PMDSEL1) );
    zan2b U287 ( .A(BUSFREE), .B(n1148), .Y(BUSFREE1) );
    zan2b U288 ( .A(RDYACK), .B(n1188), .Y(RDYACK1) );
    zan2b U289 ( .A(MADDR), .B(PCIDMA_SEL[1]), .Y(MADDR2) );
    zan2b U290 ( .A(LATCHDAT), .B(USBDMA_SEL[3]), .Y(LATCHDAT4) );
    znd2b U291 ( .A(PCIDMA_SEL[1]), .B(n1314), .Y(UGNTI2_) );
    zao2x4b U292 ( .A(MSWR4), .B(PCIDMA_SEL[3]), .C(MSWR3), .D(PCIDMA_SEL[2]), 
        .E(MSWR1), .F(n1189), .G(MSWR2), .H(PCIDMA_SEL[1]), .Y(MSWR) );
    zan2b U293 ( .A(MADDR), .B(PCIDMA_SEL[3]), .Y(MADDR4) );
    zan2b U294 ( .A(LATCHDAT), .B(USBDMA_SEL[1]), .Y(LATCHDAT2) );
    zao2x4b U295 ( .A(MRDMPLZ1), .B(n1187), .C(MRDMPLZ4), .D(PCIDMA_SEL[3]), 
        .E(MRDMPLZ2), .F(PCIDMA_SEL[1]), .G(MRDMPLZ3), .H(PCIDMA_SEL[2]), .Y(
        MRDMPLZ) );
    zan2b U296 ( .A(RDYACK), .B(PCIDMA_SEL[2]), .Y(RDYACK3) );
    zan2b U297 ( .A(LATCHDAT), .B(USBDMA_SEL[4]), .Y(LATCHDAT5) );
    zor4b U298 ( .A(BIST_ERR_S4), .B(BIST_ERR_S3), .C(BIST_ERR_S1), .D(
        BIST_ERR_S2), .Y(BIST_ERR_S) );
    zao2x4b U299 ( .A(CREQ4), .B(PCIDMA_SEL[3]), .C(CREQ1), .D(n1148), .E(
        CREQ2), .F(PCIDMA_SEL[1]), .G(CREQ3), .H(PCIDMA_SEL[2]), .Y(CREQ) );
    zan2b U300 ( .A(PMDSEL), .B(PCIDMA_SEL[3]), .Y(PMDSEL4) );
    zan2b U301 ( .A(USBDMA_SEL[1]), .B(USBPOP), .Y(USBPOP2) );
    zan2b U302 ( .A(PMDSEL), .B(PCIDMA_SEL[1]), .Y(PMDSEL2) );
    zan2b U303 ( .A(PMSTR), .B(PCIDMA_SEL[2]), .Y(PMSTR3) );
    zan2b U304 ( .A(BUSFREE), .B(PCIDMA_SEL[2]), .Y(BUSFREE3) );
    zao2x4b U305 ( .A(COMPL2), .B(PCIDMA_SEL[1]), .C(COMPL4), .D(PCIDMA_SEL[3]
        ), .E(COMPL3), .F(PCIDMA_SEL[2]), .G(COMPL1), .H(n1188), .Y(COMPL) );
    zan2b U306 ( .A(USBDMA_SEL[2]), .B(USBPOP), .Y(USBPOP3) );
    zao2x4b U307 ( .A(MRDY3_), .B(PCIDMA_SEL[2]), .C(MRDY2_), .D(PCIDMA_SEL[1]
        ), .E(MRDY1_), .F(n1188), .G(MRDY4_), .H(PCIDMA_SEL[3]), .Y(MRDY_) );
    zan2b U308 ( .A(PMSTR), .B(PCIDMA_SEL[1]), .Y(PMSTR2) );
    zan2b U309 ( .A(BUSFREE), .B(PCIDMA_SEL[3]), .Y(BUSFREE4) );
    zan2b U310 ( .A(PMDSEL), .B(PCIDMA_SEL[2]), .Y(PMDSEL3) );
    zan2b U311 ( .A(RDYACK), .B(PCIDMA_SEL[1]), .Y(RDYACK2) );
    zan2b U312 ( .A(PMSTR), .B(n1189), .Y(PMSTR1) );
    zan2b U313 ( .A(LATCHDAT), .B(n1181), .Y(LATCHDAT1) );
    zan2b U314 ( .A(n1184), .B(USBPOP), .Y(USBPOP1) );
    znd2b U315 ( .A(n1187), .B(n1314), .Y(UGNTI1_) );
    zan2b U316 ( .A(TRAN_CMD1[32]), .B(n1183), .Y(n1277) );
    zan2b U317 ( .A(TRAN_CMD1[31]), .B(n1183), .Y(n1275) );
    zan2b U318 ( .A(TRAN_CMD1[30]), .B(n1183), .Y(n1273) );
    zan2b U319 ( .A(TRAN_CMD1[29]), .B(n1183), .Y(n1271) );
    zan2b U320 ( .A(TRAN_CMD1[39]), .B(n1183), .Y(n1291) );
    zan2b U321 ( .A(TRAN_CMD1[38]), .B(n1184), .Y(n1289) );
    zan2b U322 ( .A(TRAN_CMD1[37]), .B(n1184), .Y(n1287) );
    zan2b U323 ( .A(TRAN_CMD1[36]), .B(n1181), .Y(n1285) );
    zan2b U324 ( .A(TRAN_CMD1[35]), .B(n1183), .Y(n1283) );
    zan2b U325 ( .A(TRAN_CMD1[34]), .B(n1181), .Y(n1281) );
    zan2b U326 ( .A(TRAN_CMD1[33]), .B(n1183), .Y(n1279) );
    zan2b U327 ( .A(TRAN_CMD1[6]), .B(n1182), .Y(n1225) );
    zan2b U328 ( .A(TRAN_CMD1[7]), .B(n1183), .Y(n1227) );
    zan2b U329 ( .A(TRAN_CMD1[5]), .B(n1182), .Y(n1223) );
    zan2b U330 ( .A(TRAN_CMD1[8]), .B(n1184), .Y(n1229) );
    zan2b U331 ( .A(TRAN_CMD1[9]), .B(n1181), .Y(n1231) );
    zan2b U332 ( .A(TRAN_CMD1[14]), .B(n1183), .Y(n1241) );
    zan2b U333 ( .A(TRAN_CMD1[13]), .B(n1182), .Y(n1239) );
    zan2b U334 ( .A(TRAN_CMD1[11]), .B(n1184), .Y(n1235) );
    zan2b U335 ( .A(TRAN_CMD1[10]), .B(n1182), .Y(n1233) );
    zan2b U336 ( .A(TRAN_CMD1[12]), .B(n1183), .Y(n1237) );
    zan2b U337 ( .A(TRAN_CMD5[45]), .B(n1176), .Y(n1315) );
    zan2b U338 ( .A(TRAN_CMD5[44]), .B(n1174), .Y(n1316) );
    zan2b U339 ( .A(TRAN_CMD5[42]), .B(n1174), .Y(n1317) );
    zan2b U340 ( .A(TRAN_CMD1[50]), .B(n1182), .Y(n1318) );
    zan2b U341 ( .A(TRAN_CMD5[40]), .B(n1175), .Y(n1319) );
    zan2b U342 ( .A(TRAN_CMD1[21]), .B(n1184), .Y(n1255) );
    zan2b U343 ( .A(TRAN_CMD1[20]), .B(n1181), .Y(n1253) );
    zan2b U344 ( .A(TRAN_CMD1[19]), .B(n1183), .Y(n1251) );
    zan2b U345 ( .A(TRAN_CMD1[18]), .B(n1181), .Y(n1249) );
    zan2b U346 ( .A(TRAN_CMD1[17]), .B(n1184), .Y(n1247) );
    zan2b U347 ( .A(TRAN_CMD1[16]), .B(n1182), .Y(n1245) );
    zan2b U348 ( .A(TRAN_CMD1[15]), .B(n1183), .Y(n1243) );
    zan2b U349 ( .A(TRAN_CMD1[28]), .B(n1182), .Y(n1269) );
    zan2b U350 ( .A(TRAN_CMD1[27]), .B(n1181), .Y(n1267) );
    zan2b U351 ( .A(TRAN_CMD1[26]), .B(n1181), .Y(n1265) );
    zan2b U352 ( .A(TRAN_CMD1[25]), .B(n1182), .Y(n1263) );
    zan2b U353 ( .A(TRAN_CMD1[24]), .B(n1181), .Y(n1261) );
    zan2b U354 ( .A(TRAN_CMD1[23]), .B(n1182), .Y(n1259) );
    zan2b U355 ( .A(TRAN_CMD1[22]), .B(n1181), .Y(n1257) );
    zan2b U356 ( .A(HOSTDAT1[7]), .B(n1182), .Y(n1309) );
    zan2b U357 ( .A(HOSTDAT1[6]), .B(n1181), .Y(n1307) );
    zan2b U358 ( .A(HOSTDAT1[5]), .B(n1182), .Y(n1305) );
    zan2b U359 ( .A(HOSTDAT1[4]), .B(n1183), .Y(n1303) );
    zan2b U360 ( .A(HOSTDAT1[3]), .B(n1182), .Y(n1301) );
    zan2b U361 ( .A(HOSTDAT1[2]), .B(n1181), .Y(n1299) );
    zan2b U362 ( .A(HOSTDAT1[1]), .B(n1182), .Y(n1297) );
    zan2b U363 ( .A(HOSTDAT1[0]), .B(n1184), .Y(n1295) );
    zan2b U364 ( .A(TRAN_CMD1[51]), .B(n1184), .Y(n1293) );
    zan2b U365 ( .A(TRAN_CMD1[1]), .B(n1184), .Y(n1215) );
    zan2b U366 ( .A(TRAN_CMD1[2]), .B(n1184), .Y(n1217) );
    zan2b U367 ( .A(TRAN_CMD1[3]), .B(n1184), .Y(n1219) );
    zan2b U368 ( .A(TRAN_CMD1[4]), .B(n1184), .Y(n1221) );
    zivb U369 ( .A(USBDMA_SEL[1]), .Y(n1320) );
    znr2b U370 ( .A(PCIDMA_SEL[1]), .B(n1186), .Y(n1321) );
    zor3b U371 ( .A(USBDMA_SEL[2]), .B(USBDMA_SEL[1]), .C(n1183), .Y(n1322) );
    znr2b U372 ( .A(n1178), .B(TEST_PACKET), .Y(n1198) );
    zivb U373 ( .A(TEST_PACKET), .Y(n1194) );
    zan2b U374 ( .A(TRAN_CMD1[49]), .B(n1198), .Y(TRAN_MAXLEN1[9]) );
    zan2b U375 ( .A(TRAN_CMD1[48]), .B(n1198), .Y(TRAN_MAXLEN1[8]) );
    zan2b U376 ( .A(TRAN_CMD1[47]), .B(n1198), .Y(TRAN_MAXLEN1[7]) );
    zan2b U377 ( .A(TRAN_CMD1[46]), .B(n1198), .Y(TRAN_MAXLEN1[6]) );
    zan2b U378 ( .A(TRAN_CMD1[43]), .B(n1198), .Y(TRAN_MAXLEN1[3]) );
    zan2b U379 ( .A(TRAN_CMD1[41]), .B(n1198), .Y(TRAN_MAXLEN1[1]) );
    zxo2b U380 ( .A(SLQUEUEADDR[31]), .B(add_231_carry_19), .Y(n1324) );
    zao22b U381 ( .A(TRAN_BUFPTR2[9]), .B(n1149), .C(b997_10), .D(n1177), .Y(
        DMA_BUFPTR2[9]) );
    zao22b U382 ( .A(TRAN_BUFPTR2[8]), .B(n1149), .C(b997_9), .D(n1179), .Y(
        DMA_BUFPTR2[8]) );
    zao22b U383 ( .A(TRAN_BUFPTR2[7]), .B(n1149), .C(b997_8), .D(n1179), .Y(
        DMA_BUFPTR2[7]) );
    zao22b U384 ( .A(TRAN_BUFPTR2[6]), .B(n1195), .C(b997_7), .D(n1179), .Y(
        DMA_BUFPTR2[6]) );
    zao22b U385 ( .A(TRAN_BUFPTR2[5]), .B(n1149), .C(b997_6), .D(n1177), .Y(
        DMA_BUFPTR2[5]) );
    zao22b U386 ( .A(TRAN_BUFPTR2[4]), .B(n1150), .C(b997_5), .D(n1178), .Y(
        DMA_BUFPTR2[4]) );
    zao22b U387 ( .A(TRAN_BUFPTR2[3]), .B(n1195), .C(b997_4), .D(n1177), .Y(
        DMA_BUFPTR2[3]) );
    zao22b U388 ( .A(TRAN_BUFPTR2[2]), .B(n1150), .C(b997_3), .D(n1179), .Y(
        DMA_BUFPTR2[2]) );
    zao22b U389 ( .A(TRAN_BUFPTR2[19]), .B(n1195), .C(n1324), .D(n1177), .Y(
        DMA_BUFPTR2[19]) );
    zao22b U390 ( .A(TRAN_BUFPTR2[18]), .B(n1150), .C(b997_19), .D(n1178), .Y(
        DMA_BUFPTR2[18]) );
    zao22b U391 ( .A(TRAN_BUFPTR2[17]), .B(n1195), .C(b997_18), .D(n1177), .Y(
        DMA_BUFPTR2[17]) );
    zao22b U392 ( .A(TRAN_BUFPTR2[16]), .B(n1149), .C(b997_17), .D(n1179), .Y(
        DMA_BUFPTR2[16]) );
    zao22b U393 ( .A(TRAN_BUFPTR2[15]), .B(n1195), .C(b997_16), .D(n1177), .Y(
        DMA_BUFPTR2[15]) );
    zao22b U394 ( .A(TRAN_BUFPTR2[14]), .B(n1150), .C(b997_15), .D(n1178), .Y(
        DMA_BUFPTR2[14]) );
    zao22b U395 ( .A(TRAN_BUFPTR2[13]), .B(n1149), .C(b997_14), .D(n1178), .Y(
        DMA_BUFPTR2[13]) );
    zao22b U396 ( .A(TRAN_BUFPTR2[12]), .B(n1149), .C(b997_13), .D(n1179), .Y(
        DMA_BUFPTR2[12]) );
    zao22b U397 ( .A(TRAN_BUFPTR2[11]), .B(n1149), .C(b997_12), .D(n1177), .Y(
        DMA_BUFPTR2[11]) );
    zao22b U398 ( .A(TRAN_BUFPTR2[10]), .B(n1150), .C(b997_11), .D(n1179), .Y(
        DMA_BUFPTR2[10]) );
    zao22b U399 ( .A(TRAN_BUFPTR2[1]), .B(n1149), .C(b997_2), .D(n1178), .Y(
        DMA_BUFPTR2[1]) );
    zmux21lb U400 ( .A(SLQUEUEADDR[12]), .B(n1325), .S(n1149), .Y(DMA_BUFPTR2
        [0]) );
    zao22b U401 ( .A(TRAN_BUFPTR1[9]), .B(n1149), .C(SLQUEUEADDR[9]), .D(n1179
        ), .Y(DMA_BUFPTR1[9]) );
    zao22b U402 ( .A(TRAN_BUFPTR1[8]), .B(n1149), .C(SLQUEUEADDR[8]), .D(n1177
        ), .Y(DMA_BUFPTR1[8]) );
    zao22b U403 ( .A(TRAN_BUFPTR1[7]), .B(n1149), .C(SLQUEUEADDR[7]), .D(n1179
        ), .Y(DMA_BUFPTR1[7]) );
    zao22b U404 ( .A(TRAN_BUFPTR1[6]), .B(n1149), .C(SLQUEUEADDR[6]), .D(n1177
        ), .Y(DMA_BUFPTR1[6]) );
    zao22b U405 ( .A(TRAN_BUFPTR1[5]), .B(n1150), .C(SLQUEUEADDR[5]), .D(n1179
        ), .Y(DMA_BUFPTR1[5]) );
    zao22b U406 ( .A(TRAN_BUFPTR1[4]), .B(n1149), .C(SLQUEUEADDR[4]), .D(n1177
        ), .Y(DMA_BUFPTR1[4]) );
    zao22b U407 ( .A(TRAN_BUFPTR1[31]), .B(n1150), .C(SLQUEUEADDR[31]), .D(
        n1179), .Y(DMA_BUFPTR1[31]) );
    zao22b U408 ( .A(TRAN_BUFPTR1[30]), .B(n1150), .C(SLQUEUEADDR[30]), .D(
        n1178), .Y(DMA_BUFPTR1[30]) );
    zao22b U409 ( .A(TRAN_BUFPTR1[3]), .B(n1150), .C(SLQUEUEADDR[3]), .D(n1178
        ), .Y(DMA_BUFPTR1[3]) );
    zao22b U410 ( .A(TRAN_BUFPTR1[29]), .B(n1150), .C(SLQUEUEADDR[29]), .D(
        n1177), .Y(DMA_BUFPTR1[29]) );
    zao22b U411 ( .A(TRAN_BUFPTR1[28]), .B(n1150), .C(SLQUEUEADDR[28]), .D(
        n1178), .Y(DMA_BUFPTR1[28]) );
    zao22b U412 ( .A(TRAN_BUFPTR1[27]), .B(n1150), .C(SLQUEUEADDR[27]), .D(
        n1177), .Y(DMA_BUFPTR1[27]) );
    zao22b U413 ( .A(TRAN_BUFPTR1[26]), .B(n1195), .C(SLQUEUEADDR[26]), .D(
        n1178), .Y(DMA_BUFPTR1[26]) );
    zao22b U414 ( .A(TRAN_BUFPTR1[25]), .B(n1150), .C(SLQUEUEADDR[25]), .D(
        n1177), .Y(DMA_BUFPTR1[25]) );
    zao22b U415 ( .A(TRAN_BUFPTR1[24]), .B(n1149), .C(SLQUEUEADDR[24]), .D(
        n1177), .Y(DMA_BUFPTR1[24]) );
    zao22b U416 ( .A(TRAN_BUFPTR1[23]), .B(n1195), .C(SLQUEUEADDR[23]), .D(
        n1177), .Y(DMA_BUFPTR1[23]) );
    zao22b U417 ( .A(TRAN_BUFPTR1[22]), .B(n1149), .C(SLQUEUEADDR[22]), .D(
        n1177), .Y(DMA_BUFPTR1[22]) );
    zao22b U418 ( .A(TRAN_BUFPTR1[21]), .B(n1195), .C(SLQUEUEADDR[21]), .D(
        n1177), .Y(DMA_BUFPTR1[21]) );
    zao22b U419 ( .A(TRAN_BUFPTR1[20]), .B(n1150), .C(SLQUEUEADDR[20]), .D(
        n1177), .Y(DMA_BUFPTR1[20]) );
    zao22b U420 ( .A(TRAN_BUFPTR1[2]), .B(n1150), .C(SLQUEUEADDR[2]), .D(n1178
        ), .Y(DMA_BUFPTR1[2]) );
    zao22b U421 ( .A(TRAN_BUFPTR1[19]), .B(n1149), .C(SLQUEUEADDR[19]), .D(
        n1177), .Y(DMA_BUFPTR1[19]) );
    zao22b U422 ( .A(TRAN_BUFPTR1[18]), .B(n1195), .C(SLQUEUEADDR[18]), .D(
        n1178), .Y(DMA_BUFPTR1[18]) );
    zao22b U423 ( .A(TRAN_BUFPTR1[17]), .B(n1150), .C(SLQUEUEADDR[17]), .D(
        n1178), .Y(DMA_BUFPTR1[17]) );
    zao22b U424 ( .A(TRAN_BUFPTR1[16]), .B(n1195), .C(SLQUEUEADDR[16]), .D(
        n1178), .Y(DMA_BUFPTR1[16]) );
    zao22b U425 ( .A(TRAN_BUFPTR1[15]), .B(n1195), .C(SLQUEUEADDR[15]), .D(
        n1179), .Y(DMA_BUFPTR1[15]) );
    zao22b U426 ( .A(TRAN_BUFPTR1[14]), .B(n1195), .C(SLQUEUEADDR[14]), .D(
        n1179), .Y(DMA_BUFPTR1[14]) );
    zao22b U427 ( .A(TRAN_BUFPTR1[13]), .B(n1195), .C(SLQUEUEADDR[13]), .D(
        n1179), .Y(DMA_BUFPTR1[13]) );
    zao22b U428 ( .A(TRAN_BUFPTR1[12]), .B(n1195), .C(SLQUEUEADDR[12]), .D(
        n1179), .Y(DMA_BUFPTR1[12]) );
    zao22b U429 ( .A(TRAN_BUFPTR1[11]), .B(n1195), .C(SLQUEUEADDR[11]), .D(
        n1179), .Y(DMA_BUFPTR1[11]) );
    zao22b U430 ( .A(TRAN_BUFPTR1[10]), .B(n1149), .C(SLQUEUEADDR[10]), .D(
        n1179), .Y(DMA_BUFPTR1[10]) );
    zao22b U431 ( .A(TRAN_BUFPTR1[1]), .B(n1149), .C(SLQUEUEADDR[1]), .D(n1179
        ), .Y(DMA_BUFPTR1[1]) );
    zao22b U432 ( .A(TRAN_BUFPTR1[0]), .B(n1195), .C(SLQUEUEADDR[0]), .D(n1179
        ), .Y(DMA_BUFPTR1[0]) );
    zao222b U433 ( .A(TRAN_CMD5[32]), .B(n1174), .C(TRAN_CMD2[32]), .D(n1193), 
        .E(TRAN_CMD4[32]), .F(n1151), .Y(n1278) );
    zao222b U434 ( .A(TRAN_CMD5[31]), .B(n1175), .C(TRAN_CMD2[31]), .D(n1191), 
        .E(TRAN_CMD4[31]), .F(n1151), .Y(n1276) );
    zao222b U435 ( .A(TRAN_CMD5[30]), .B(n1176), .C(TRAN_CMD2[30]), .D(n1193), 
        .E(TRAN_CMD4[30]), .F(n1151), .Y(n1274) );
    zao222b U436 ( .A(TRAN_CMD5[29]), .B(n1174), .C(TRAN_CMD2[29]), .D(n1192), 
        .E(TRAN_CMD4[29]), .F(n1151), .Y(n1272) );
    zao222b U437 ( .A(TRAN_CMD5[39]), .B(n1175), .C(TRAN_CMD2[39]), .D(n1193), 
        .E(TRAN_CMD4[39]), .F(n1151), .Y(n1292) );
    zao222b U438 ( .A(TRAN_CMD5[38]), .B(n1175), .C(TRAN_CMD2[38]), .D(n1193), 
        .E(TRAN_CMD4[38]), .F(n1151), .Y(n1290) );
    zao222b U439 ( .A(TRAN_CMD5[37]), .B(n1175), .C(TRAN_CMD2[37]), .D(n1192), 
        .E(TRAN_CMD4[37]), .F(n1151), .Y(n1288) );
    zao222b U440 ( .A(TRAN_CMD5[36]), .B(n1174), .C(TRAN_CMD2[36]), .D(n1192), 
        .E(TRAN_CMD4[36]), .F(n1151), .Y(n1286) );
    zao222b U441 ( .A(TRAN_CMD5[35]), .B(n1176), .C(TRAN_CMD2[35]), .D(n1191), 
        .E(TRAN_CMD4[35]), .F(n1151), .Y(n1284) );
    zao222b U442 ( .A(TRAN_CMD5[34]), .B(n1176), .C(TRAN_CMD2[34]), .D(n1192), 
        .E(TRAN_CMD4[34]), .F(n1151), .Y(n1282) );
    zao222b U443 ( .A(TRAN_CMD5[33]), .B(n1176), .C(TRAN_CMD2[33]), .D(n1191), 
        .E(TRAN_CMD4[33]), .F(n1151), .Y(n1280) );
    zao222b U444 ( .A(TRAN_CMD5[6]), .B(n1174), .C(TRAN_CMD2[6]), .D(n1193), 
        .E(TRAN_CMD4[6]), .F(n1151), .Y(n1226) );
    zao222b U445 ( .A(TRAN_CMD5[7]), .B(n1174), .C(TRAN_CMD2[7]), .D(n1191), 
        .E(TRAN_CMD4[7]), .F(n1151), .Y(n1228) );
    zao222b U446 ( .A(TRAN_CMD5[5]), .B(n1176), .C(TRAN_CMD2[5]), .D(n1191), 
        .E(TRAN_CMD4[5]), .F(n1151), .Y(n1224) );
    zao222b U447 ( .A(TRAN_CMD5[8]), .B(n1174), .C(TRAN_CMD2[8]), .D(n1193), 
        .E(TRAN_CMD4[8]), .F(n1153), .Y(n1230) );
    zao222b U448 ( .A(TRAN_CMD5[9]), .B(n1175), .C(TRAN_CMD2[9]), .D(n1191), 
        .E(TRAN_CMD4[9]), .F(n1151), .Y(n1232) );
    zao222b U449 ( .A(TRAN_CMD5[14]), .B(n1175), .C(TRAN_CMD2[14]), .D(n1193), 
        .E(TRAN_CMD4[14]), .F(n1151), .Y(n1242) );
    zao222b U450 ( .A(TRAN_CMD5[13]), .B(n1176), .C(TRAN_CMD2[13]), .D(n1192), 
        .E(TRAN_CMD4[13]), .F(n1151), .Y(n1240) );
    zao222b U451 ( .A(TRAN_CMD5[11]), .B(n1174), .C(TRAN_CMD2[11]), .D(n1193), 
        .E(TRAN_CMD4[11]), .F(n1151), .Y(n1236) );
    zao222b U452 ( .A(TRAN_CMD5[10]), .B(n1175), .C(TRAN_CMD2[10]), .D(n1193), 
        .E(TRAN_CMD4[10]), .F(n1151), .Y(n1234) );
    zao222b U453 ( .A(TRAN_CMD5[12]), .B(n1176), .C(TRAN_CMD2[12]), .D(n1191), 
        .E(TRAN_CMD4[12]), .F(n1152), .Y(n1238) );
    zao211b U454 ( .A(TRAN_CMD2[45]), .B(n1193), .C(TEST_PACKET), .D(n1315), 
        .Y(n1203) );
    zao222b U455 ( .A(TRAN_CMD3[45]), .B(n1157), .C(TRAN_CMD4[45]), .D(n1152), 
        .E(TRAN_CMD1[45]), .F(n1184), .Y(n1204) );
    zao211b U456 ( .A(TRAN_CMD2[44]), .B(n1191), .C(TEST_PACKET), .D(n1316), 
        .Y(n1205) );
    zao222b U457 ( .A(TRAN_CMD3[44]), .B(n1156), .C(TRAN_CMD4[44]), .D(n1152), 
        .E(TRAN_CMD1[44]), .F(n1181), .Y(n1206) );
    zao211b U458 ( .A(TRAN_CMD2[42]), .B(n1192), .C(TEST_PACKET), .D(n1317), 
        .Y(n1208) );
    zao222b U459 ( .A(TRAN_CMD3[42]), .B(n1155), .C(TRAN_CMD4[42]), .D(n1152), 
        .E(TRAN_CMD1[42]), .F(n1184), .Y(n1209) );
    zao222b U460 ( .A(TRAN_CMD5[50]), .B(n1175), .C(TRAN_CMD2[50]), .D(n1191), 
        .E(TRAN_CMD4[50]), .F(n1152), .Y(n1326) );
    zao211b U461 ( .A(TRAN_CMD2[40]), .B(n1191), .C(TEST_PACKET), .D(n1319), 
        .Y(n1211) );
    zao222b U462 ( .A(TRAN_CMD3[40]), .B(n1157), .C(TRAN_CMD4[40]), .D(n1152), 
        .E(TRAN_CMD1[40]), .F(n1181), .Y(n1212) );
    zao222b U463 ( .A(TRAN_CMD5[0]), .B(n1176), .C(TRAN_CMD2[0]), .D(n1192), 
        .E(TRAN_CMD4[0]), .F(n1153), .Y(n1311) );
    zao22b U464 ( .A(TRAN_CMD1[0]), .B(n1182), .C(TRAN_CMD3[0]), .D(n1155), 
        .Y(n1312) );
    zao222b U465 ( .A(TRAN_CMD5[21]), .B(n1175), .C(TRAN_CMD2[21]), .D(n1193), 
        .E(TRAN_CMD4[21]), .F(n1153), .Y(n1256) );
    zao222b U466 ( .A(TRAN_CMD5[20]), .B(n1174), .C(TRAN_CMD2[20]), .D(n1192), 
        .E(TRAN_CMD4[20]), .F(n1153), .Y(n1254) );
    zao222b U467 ( .A(TRAN_CMD5[19]), .B(n1174), .C(TRAN_CMD2[19]), .D(n1193), 
        .E(TRAN_CMD4[19]), .F(n1153), .Y(n1252) );
    zao222b U468 ( .A(TRAN_CMD5[18]), .B(n1176), .C(TRAN_CMD2[18]), .D(n1191), 
        .E(TRAN_CMD4[18]), .F(n1152), .Y(n1250) );
    zao222b U469 ( .A(TRAN_CMD5[17]), .B(n1174), .C(TRAN_CMD2[17]), .D(n1192), 
        .E(TRAN_CMD4[17]), .F(n1153), .Y(n1248) );
    zao222b U470 ( .A(TRAN_CMD5[16]), .B(n1174), .C(TRAN_CMD2[16]), .D(n1192), 
        .E(TRAN_CMD4[16]), .F(n1153), .Y(n1246) );
    zao222b U471 ( .A(TRAN_CMD5[15]), .B(n1176), .C(TRAN_CMD2[15]), .D(n1191), 
        .E(TRAN_CMD4[15]), .F(n1153), .Y(n1244) );
    zao222b U472 ( .A(TRAN_CMD5[28]), .B(n1175), .C(TRAN_CMD2[28]), .D(n1192), 
        .E(TRAN_CMD4[28]), .F(n1153), .Y(n1270) );
    zao222b U473 ( .A(TRAN_CMD5[27]), .B(n1174), .C(TRAN_CMD2[27]), .D(n1193), 
        .E(TRAN_CMD4[27]), .F(n1153), .Y(n1268) );
    zao222b U474 ( .A(TRAN_CMD5[26]), .B(n1175), .C(TRAN_CMD2[26]), .D(n1191), 
        .E(TRAN_CMD4[26]), .F(n1153), .Y(n1266) );
    zao222b U475 ( .A(TRAN_CMD5[25]), .B(n1175), .C(TRAN_CMD2[25]), .D(n1191), 
        .E(TRAN_CMD4[25]), .F(n1153), .Y(n1264) );
    zao222b U476 ( .A(TRAN_CMD5[24]), .B(n1175), .C(TRAN_CMD2[24]), .D(n1193), 
        .E(TRAN_CMD4[24]), .F(n1153), .Y(n1262) );
    zao222b U477 ( .A(TRAN_CMD5[23]), .B(n1175), .C(TRAN_CMD2[23]), .D(n1192), 
        .E(TRAN_CMD4[23]), .F(n1153), .Y(n1260) );
    zao222b U478 ( .A(TRAN_CMD5[22]), .B(n1176), .C(TRAN_CMD2[22]), .D(n1192), 
        .E(TRAN_CMD4[22]), .F(n1153), .Y(n1258) );
    zao222b U479 ( .A(HOSTDAT5[7]), .B(n1174), .C(HOSTDAT2[7]), .D(n1191), .E(
        HOSTDAT4[7]), .F(n1153), .Y(n1310) );
    zao222b U480 ( .A(HOSTDAT5[6]), .B(n1175), .C(HOSTDAT2[6]), .D(n1192), .E(
        HOSTDAT4[6]), .F(n1152), .Y(n1308) );
    zao222b U481 ( .A(HOSTDAT5[5]), .B(n1175), .C(HOSTDAT2[5]), .D(n1193), .E(
        HOSTDAT4[5]), .F(n1153), .Y(n1306) );
    zao222b U482 ( .A(HOSTDAT5[4]), .B(n1176), .C(HOSTDAT2[4]), .D(n1191), .E(
        HOSTDAT4[4]), .F(n1152), .Y(n1304) );
    zao222b U483 ( .A(HOSTDAT5[3]), .B(n1174), .C(HOSTDAT2[3]), .D(n1192), .E(
        HOSTDAT4[3]), .F(n1153), .Y(n1302) );
    zao222b U484 ( .A(HOSTDAT5[2]), .B(n1176), .C(HOSTDAT2[2]), .D(n1193), .E(
        HOSTDAT4[2]), .F(n1152), .Y(n1300) );
    zao222b U485 ( .A(HOSTDAT5[1]), .B(n1174), .C(HOSTDAT2[1]), .D(n1191), .E(
        HOSTDAT4[1]), .F(n1153), .Y(n1298) );
    zao222b U486 ( .A(HOSTDAT5[0]), .B(n1176), .C(HOSTDAT2[0]), .D(n1192), .E(
        HOSTDAT4[0]), .F(n1152), .Y(n1296) );
    zao222b U487 ( .A(TRAN_CMD5[51]), .B(n1176), .C(TRAN_CMD2[51]), .D(n1193), 
        .E(TRAN_CMD4[51]), .F(n1152), .Y(n1294) );
    zao222b U488 ( .A(TRAN_CMD5[1]), .B(n1175), .C(TRAN_CMD2[1]), .D(n1191), 
        .E(TRAN_CMD4[1]), .F(n1152), .Y(n1216) );
    zao222b U489 ( .A(TRAN_CMD5[2]), .B(n1176), .C(TRAN_CMD2[2]), .D(n1193), 
        .E(TRAN_CMD4[2]), .F(n1152), .Y(n1218) );
    zao222b U490 ( .A(TRAN_CMD5[3]), .B(n1176), .C(TRAN_CMD2[3]), .D(n1192), 
        .E(TRAN_CMD4[3]), .F(n1153), .Y(n1220) );
    zao222b U491 ( .A(TRAN_CMD5[4]), .B(n1174), .C(TRAN_CMD2[4]), .D(n1192), 
        .E(TRAN_CMD4[4]), .F(n1151), .Y(n1222) );
    zivb U492 ( .A(UGNTI_), .Y(n1314) );
    zivb U493 ( .A(SLAVE_ACT), .Y(n1313) );
    znr2b U494 ( .A(n1178), .B(n1194), .Y(n1196) );
    zao2x4b U495 ( .A(TRAN_CMD3[49]), .B(n1157), .C(TRAN_CMD4[49]), .D(n1152), 
        .E(TRAN_CMD5[49]), .F(n1176), .G(TRAN_CMD2[49]), .H(n1193), .Y(n1199)
         );
    zao2x4b U496 ( .A(TRAN_CMD3[48]), .B(n1155), .C(TRAN_CMD4[48]), .D(n1152), 
        .E(TRAN_CMD5[48]), .F(n1175), .G(TRAN_CMD2[48]), .H(n1193), .Y(n1200)
         );
    zao2x4b U497 ( .A(TRAN_CMD3[47]), .B(n1156), .C(TRAN_CMD4[47]), .D(n1152), 
        .E(TRAN_CMD5[47]), .F(n1174), .G(TRAN_CMD2[47]), .H(n1192), .Y(n1201)
         );
    zao2x4b U498 ( .A(TRAN_CMD3[46]), .B(n1157), .C(TRAN_CMD4[46]), .D(n1152), 
        .E(TRAN_CMD5[46]), .F(n1175), .G(TRAN_CMD2[46]), .H(n1192), .Y(n1202)
         );
    zao2x4b U499 ( .A(TRAN_CMD3[43]), .B(n1156), .C(TRAN_CMD4[43]), .D(n1152), 
        .E(TRAN_CMD5[43]), .F(n1176), .G(TRAN_CMD2[43]), .H(n1191), .Y(n1207)
         );
    zao211b U500 ( .A(TRAN_CMD3[50]), .B(n1157), .C(n1318), .D(n1326), .Y(
        n1197) );
    zao2x4b U501 ( .A(TRAN_CMD3[41]), .B(n1155), .C(TRAN_CMD4[41]), .D(n1152), 
        .E(TRAN_CMD5[41]), .F(n1174), .G(TRAN_CMD2[41]), .H(n1191), .Y(n1210)
         );
    zivb U502 ( .A(TRAN_BUFPTR2[0]), .Y(n1325) );
endmodule


module HS_CLKCTL ( RUN, EHCI_IDLE, USBDMA_SEL, SLAVEMODE, TEST_EYE_EN, 
    PTstCtrl_A_3, PTstCtrl_A_2, PTstCtrl_A_1, PTstCtrl_A_0, PTstCtrl_B_3, 
    PTstCtrl_B_2, PTstCtrl_B_1, PTstCtrl_B_0, PTstCtrl_C_3, PTstCtrl_C_2, 
    PTstCtrl_C_1, PTstCtrl_C_0, PTstCtrl_D_3, PTstCtrl_D_2, PTstCtrl_D_1, 
    PTstCtrl_D_0, PTstCtrl_E_3, PTstCtrl_E_2, PTstCtrl_E_1, PTstCtrl_E_0, 
    PTstCtrl_F_3, PTstCtrl_F_2, PTstCtrl_F_1, PTstCtrl_F_0, PTstCtrl_G_3, 
    PTstCtrl_G_2, PTstCtrl_G_1, PTstCtrl_G_0, PTstCtrl_H_3, PTstCtrl_H_2, 
    PTstCtrl_H_1, PTstCtrl_H_0, HCIREQ1, HCIREQ2, SLHCIREQ, BIST_RUN, UADS, 
    TD_PARSE_GO1, TD_PARSE_GO2, TD_PARSE_GO3, TD_PARSE_GO4, TD_IDLE1, TD_IDLE2, 
    TD_IDLE3, TD_IDLE4, EHCIFLOW_PCLK_EN, MAC_CLK60M_EN, EHCI_DMA_EN1, 
    EHCI_DMA_EN2, EHCI_DMA_EN3, EHCI_DMA_EN4, DMA_CLK60M_EN1, DMA_CLK60M_EN2, 
    DMA_CLK60M_EN3, DMA_CLK60M_EN4, DMA_IDLE1, DMA_IDLE2, DMA_IDLE3, DMA_IDLE4, 
    PCIS_ACT, PCLK33_EN, TX_PERIOD, ASKREPLY, HS_MAC_TX_EN, HS_MAC_RX_EN, 
    AUTOCHK, AUTOCHK_CLK60M_EN, EN_DBG_PORT, DBG_OWNER, DBG_ENABLE, DBG_GO, 
    DBG_IDLE, DBG_PCLK_EN, DBG_CLK60M_EN, CLKOFF_EN, PCLK66, PCLK33, CLK60M, 
    HRST_, ATPG_ENI );
input  [4:0] USBDMA_SEL;
input  RUN, EHCI_IDLE, SLAVEMODE, TEST_EYE_EN, PTstCtrl_A_3, PTstCtrl_A_2, 
    PTstCtrl_A_1, PTstCtrl_A_0, PTstCtrl_B_3, PTstCtrl_B_2, PTstCtrl_B_1, 
    PTstCtrl_B_0, PTstCtrl_C_3, PTstCtrl_C_2, PTstCtrl_C_1, PTstCtrl_C_0, 
    PTstCtrl_D_3, PTstCtrl_D_2, PTstCtrl_D_1, PTstCtrl_D_0, PTstCtrl_E_3, 
    PTstCtrl_E_2, PTstCtrl_E_1, PTstCtrl_E_0, PTstCtrl_F_3, PTstCtrl_F_2, 
    PTstCtrl_F_1, PTstCtrl_F_0, PTstCtrl_G_3, PTstCtrl_G_2, PTstCtrl_G_1, 
    PTstCtrl_G_0, PTstCtrl_H_3, PTstCtrl_H_2, PTstCtrl_H_1, PTstCtrl_H_0, 
    HCIREQ1, HCIREQ2, SLHCIREQ, BIST_RUN, UADS, TD_PARSE_GO1, TD_PARSE_GO2, 
    TD_PARSE_GO3, TD_PARSE_GO4, TD_IDLE1, TD_IDLE2, TD_IDLE3, TD_IDLE4, 
    DMA_IDLE1, DMA_IDLE2, DMA_IDLE3, DMA_IDLE4, PCIS_ACT, TX_PERIOD, ASKREPLY, 
    AUTOCHK, EN_DBG_PORT, DBG_OWNER, DBG_ENABLE, DBG_GO, DBG_IDLE, CLKOFF_EN, 
    PCLK66, PCLK33, CLK60M, HRST_, ATPG_ENI;
output EHCIFLOW_PCLK_EN, MAC_CLK60M_EN, EHCI_DMA_EN1, EHCI_DMA_EN2, 
    EHCI_DMA_EN3, EHCI_DMA_EN4, DMA_CLK60M_EN1, DMA_CLK60M_EN2, DMA_CLK60M_EN3, 
    DMA_CLK60M_EN4, PCLK33_EN, HS_MAC_TX_EN, HS_MAC_RX_EN, AUTOCHK_CLK60M_EN, 
    DBG_PCLK_EN, DBG_CLK60M_EN;
    wire SPAREO6, UADS_T, DMA_CLK60M_EN4_P1189, PCLK33_EN_2T, EHCI_DMA_EN1_P, 
        HS_MAC_RX_EN_P771, DBG_PCLK_EN_P, MAC_CLK60M_EN_P, TEST_FORCE_ENABLE, 
        UADS_EN, SPAREO0_, SPAREO8, TEST_SE0_NAK, HS_MAC_TX_EN_2T, 
        HS_MAC_RX_EN_T, DMA_CLK60M_EN3_P, EHCI_DMA_EN2_2T, SPAREO1, 
        DMA_CLK60M_EN2_P, HS_MAC_TX_EN_T, SPAREO9, EHCI_DMA_EN4_P, 
        EHCIFLOW_PCLK_EN_T, PCLK33_EN_T1267, EHCI_DMA_EN3_2T, 
        EHCIFLOW_PCLK_EN_P501, SPAREO0, UADS_2T, EHCI_DMA_EN3_T, 
        DBG_PCLK_EN_P1321, SPAREO7, EHCI_DMA_EN2_T, EHCI_DMA_EN2_P875, 
        DMA_CLK60M_EN2_P1177, HS_MAC_RX_EN_2T, SPAREO5, DMA_CLK60M_EN1_P1171, 
        DBG_CLK60M_EN_P, HS_MAC_RX_EN_P, DBG_PCLK_EN_T, MAC_CLK60M_EN_T, 
        DMA_CLK60M_EN4_P, EHCI_DMA_EN1_T, DBG_PCLK_EN_2T, EHCI_DMA_EN4_P887, 
        SPAREO2, TEST_K, MAC_CLK60M_EN_2T, TEST_J, EHCI_DMA_EN1_P869, SPAREO3, 
        EHCI_DMA_EN2_P, DBG_CLK60M_EN_P1413, SPAREO1_, EHCI_DMA_EN3_P881, 
        EHCI_DMA_EN3_P, PCLK33_EN_T, EHCI_DMA_EN4_2T, HS_MAC_TX_EN_P701, 
        PCLK33_EN_3T, SPAREO4, MAC_CLK60M_EN_P593, EHCIFLOW_PCLK_EN_2T, 
        DMA_CLK60M_EN1_P, EHCIFLOW_PCLK_EN_P, DMA_CLK60M_EN3_P1183, 
        AUTOCHK_CLK60M_EN_P, EHCI_DMA_EN4_T, HS_MAC_TX_EN_P, EHCI_DMA_EN1_2T, 
        n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, 
        n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, 
        n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521;
    zivb SPARE887 ( .A(SPAREO4), .Y(SPAREO5) );
    zdffrb SPARE880 ( .CK(PCLK66), .D(1'b0), .R(HRST_), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE889 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zdffrb SPARE881 ( .CK(CLK60M), .D(SPAREO7), .R(HRST_), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zivb SPARE888 ( .A(SPAREO5), .Y(SPAREO6) );
    znr3b SPARE886 ( .A(SPAREO2), .B(UADS_EN), .C(SPAREO0_), .Y(SPAREO4) );
    zoai21b SPARE884 ( .A(SPAREO0), .B(SPAREO8), .C(TEST_K), .Y(SPAREO9) );
    zaoi211b SPARE883 ( .A(SPAREO4), .B(1'b0), .C(SPAREO6), .D(TEST_J), .Y(
        SPAREO8) );
    zaoi211b SPARE882 ( .A(SPAREO0), .B(TEST_EYE_EN), .C(SPAREO1_), .D(
        TEST_SE0_NAK), .Y(SPAREO2) );
    zoai21b SPARE885 ( .A(SPAREO1), .B(TEST_FORCE_ENABLE), .C(SPAREO9), .Y(
        SPAREO3) );
    zdffqrb_ AUTOCHK_CLK60M_EN_P_reg ( .CK(CLK60M), .D(AUTOCHK), .R(HRST_), 
        .Q(AUTOCHK_CLK60M_EN_P) );
    zdffqrb_ PCLK33_EN_3T_reg ( .CK(PCLK33), .D(PCLK33_EN_2T), .R(HRST_), .Q(
        PCLK33_EN_3T) );
    zdffqrb_ UADS_2T_reg ( .CK(PCLK66), .D(UADS_T), .R(HRST_), .Q(UADS_2T) );
    zdffqrb_ PCLK33_EN_2T_reg ( .CK(PCLK33), .D(PCLK33_EN_T), .R(HRST_), .Q(
        PCLK33_EN_2T) );
    zdffqrb_ UADS_T_reg ( .CK(PCLK66), .D(UADS), .R(HRST_), .Q(UADS_T) );
    zdffqrb_ PCLK33_EN_T_reg ( .CK(PCLK33), .D(PCLK33_EN_T1267), .R(HRST_), 
        .Q(PCLK33_EN_T) );
    zdffqrb_ DBG_CLK60M_EN_P_reg ( .CK(CLK60M), .D(DBG_CLK60M_EN_P1413), .R(
        HRST_), .Q(DBG_CLK60M_EN_P) );
    zor5b U377 ( .A(ATPG_ENI), .B(PCLK33_EN_3T), .C(PCIS_ACT), .D(PCLK33_EN_T), 
        .E(PCLK33_EN_2T), .Y(PCLK33_EN) );
    zor2b U378 ( .A(ATPG_ENI), .B(n1492), .Y(EHCI_DMA_EN1) );
    zor2b U379 ( .A(TX_PERIOD), .B(n1493), .Y(HS_MAC_TX_EN_P701) );
    zor4b U380 ( .A(DBG_PCLK_EN_P), .B(DBG_PCLK_EN_T), .C(ATPG_ENI), .D(
        DBG_PCLK_EN_2T), .Y(DBG_PCLK_EN) );
    zor5b U381 ( .A(ATPG_ENI), .B(HS_MAC_RX_EN_2T), .C(HS_MAC_RX_EN_P), .D(
        HS_MAC_RX_EN_T), .E(n1493), .Y(HS_MAC_RX_EN) );
    zor3b U382 ( .A(UADS_2T), .B(UADS), .C(UADS_T), .Y(UADS_EN) );
    zor5b U383 ( .A(ATPG_ENI), .B(HS_MAC_TX_EN_P701), .C(HS_MAC_TX_EN_2T), .D(
        HS_MAC_TX_EN_T), .E(HS_MAC_TX_EN_P), .Y(HS_MAC_TX_EN) );
    zor4b U384 ( .A(USBDMA_SEL[4]), .B(DBG_PCLK_EN_P1321), .C(DBG_PCLK_EN), 
        .D(AUTOCHK), .Y(DBG_CLK60M_EN_P1413) );
    zor3b U385 ( .A(USBDMA_SEL[2]), .B(n1493), .C(n1494), .Y(
        DMA_CLK60M_EN3_P1183) );
    zor2b U386 ( .A(DMA_CLK60M_EN4_P), .B(ATPG_ENI), .Y(DMA_CLK60M_EN4) );
    zor3b U387 ( .A(USBDMA_SEL[0]), .B(n1493), .C(n1492), .Y(
        DMA_CLK60M_EN1_P1171) );
    zor4b U388 ( .A(MAC_CLK60M_EN_P), .B(MAC_CLK60M_EN_T), .C(ATPG_ENI), .D(
        MAC_CLK60M_EN_2T), .Y(MAC_CLK60M_EN) );
    zor2b U389 ( .A(DBG_CLK60M_EN_P), .B(ATPG_ENI), .Y(DBG_CLK60M_EN) );
    zor4b U390 ( .A(EHCIFLOW_PCLK_EN_P), .B(EHCIFLOW_PCLK_EN_T), .C(ATPG_ENI), 
        .D(EHCIFLOW_PCLK_EN_2T), .Y(EHCIFLOW_PCLK_EN) );
    zor5b U391 ( .A(HCIREQ1), .B(TD_PARSE_GO1), .C(n1495), .D(SLHCIREQ), .E(
        n1496), .Y(EHCI_DMA_EN1_P869) );
    zan2b U392 ( .A(n1497), .B(n1498), .Y(TEST_SE0_NAK) );
    zor3b U393 ( .A(TD_PARSE_GO4), .B(n1499), .C(n1500), .Y(EHCI_DMA_EN4_P887)
         );
    zor3b U394 ( .A(TD_PARSE_GO2), .B(n1499), .C(n1501), .Y(EHCI_DMA_EN2_P875)
         );
    zao211b U395 ( .A(EN_DBG_PORT), .B(n1502), .C(UADS_EN), .D(n1493), .Y(
        DBG_PCLK_EN_P1321) );
    zor2b U396 ( .A(DMA_CLK60M_EN1_P), .B(ATPG_ENI), .Y(DMA_CLK60M_EN1) );
    zor3b U397 ( .A(AUTOCHK), .B(ASKREPLY), .C(n1493), .Y(HS_MAC_RX_EN_P771)
         );
    zor2b U398 ( .A(ATPG_ENI), .B(n1503), .Y(EHCI_DMA_EN2) );
    zor2b U399 ( .A(DMA_CLK60M_EN3_P), .B(ATPG_ENI), .Y(DMA_CLK60M_EN3) );
    zor2b U400 ( .A(n1504), .B(UADS), .Y(EHCIFLOW_PCLK_EN_P501) );
    zor2b U401 ( .A(n1493), .B(PCIS_ACT), .Y(PCLK33_EN_T1267) );
    zor3b U402 ( .A(USBDMA_SEL[1]), .B(n1493), .C(n1503), .Y(
        DMA_CLK60M_EN2_P1177) );
    zor4b U403 ( .A(TEST_J), .B(n1504), .C(TEST_K), .D(TEST_EYE_EN), .Y(
        MAC_CLK60M_EN_P593) );
    zor2b U404 ( .A(ATPG_ENI), .B(n1505), .Y(EHCI_DMA_EN4) );
    zor3b U405 ( .A(ATPG_ENI), .B(AUTOCHK_CLK60M_EN_P), .C(n1493), .Y(
        AUTOCHK_CLK60M_EN) );
    zor2b U406 ( .A(DMA_CLK60M_EN2_P), .B(ATPG_ENI), .Y(DMA_CLK60M_EN2) );
    zor3b U407 ( .A(USBDMA_SEL[3]), .B(n1493), .C(n1505), .Y(
        DMA_CLK60M_EN4_P1189) );
    zor4b U408 ( .A(TD_PARSE_GO3), .B(HCIREQ2), .C(n1499), .D(n1506), .Y(
        EHCI_DMA_EN3_P881) );
    zor2b U409 ( .A(ATPG_ENI), .B(n1494), .Y(EHCI_DMA_EN3) );
    zan3b U410 ( .A(DBG_OWNER), .B(DBG_ENABLE), .C(EN_DBG_PORT), .Y(n1507) );
    zor5b U411 ( .A(PTstCtrl_H_2), .B(PTstCtrl_G_2), .C(PTstCtrl_F_2), .D(
        PTstCtrl_C_2), .E(n1509), .Y(n1508) );
    zor5b U412 ( .A(PTstCtrl_D_3), .B(PTstCtrl_G_3), .C(PTstCtrl_F_3), .D(
        PTstCtrl_E_3), .E(n1511), .Y(n1510) );
    zan3b U413 ( .A(n1512), .B(n1513), .C(n1514), .Y(n1497) );
    zor5b U414 ( .A(PTstCtrl_B_0), .B(PTstCtrl_H_0), .C(PTstCtrl_G_0), .D(
        PTstCtrl_A_0), .E(n1515), .Y(n1498) );
    zor5b U415 ( .A(PTstCtrl_H_1), .B(PTstCtrl_C_1), .C(PTstCtrl_A_1), .D(
        PTstCtrl_B_1), .E(n1516), .Y(n1512) );
    zor2b U416 ( .A(n1512), .B(n1510), .Y(n1517) );
    zivb U417 ( .A(CLKOFF_EN), .Y(n1493) );
    zivb U418 ( .A(EHCI_IDLE), .Y(n1518) );
    zor4b U419 ( .A(n1507), .B(n1493), .C(n1518), .D(n1519), .Y(n1504) );
    zor3b U420 ( .A(UADS_EN), .B(BIST_RUN), .C(n1493), .Y(n1499) );
    zor3b U421 ( .A(EHCI_DMA_EN4_2T), .B(EHCI_DMA_EN4_P), .C(EHCI_DMA_EN4_T), 
        .Y(n1505) );
    zor3b U422 ( .A(EHCI_DMA_EN3_P), .B(EHCI_DMA_EN3_T), .C(EHCI_DMA_EN3_2T), 
        .Y(n1494) );
    zor3b U423 ( .A(EHCI_DMA_EN2_P), .B(EHCI_DMA_EN2_T), .C(EHCI_DMA_EN2_2T), 
        .Y(n1503) );
    zor3b U424 ( .A(EHCI_DMA_EN1_P), .B(EHCI_DMA_EN1_T), .C(EHCI_DMA_EN1_2T), 
        .Y(n1492) );
    zor4b U425 ( .A(PTstCtrl_D_0), .B(PTstCtrl_E_0), .C(PTstCtrl_F_0), .D(
        PTstCtrl_C_0), .Y(n1515) );
    zor4b U426 ( .A(PTstCtrl_D_1), .B(PTstCtrl_F_1), .C(PTstCtrl_G_1), .D(
        PTstCtrl_E_1), .Y(n1516) );
    zor4b U427 ( .A(PTstCtrl_B_2), .B(PTstCtrl_D_2), .C(PTstCtrl_E_2), .D(
        PTstCtrl_A_2), .Y(n1509) );
    zor4b U428 ( .A(PTstCtrl_A_3), .B(PTstCtrl_B_3), .C(PTstCtrl_H_3), .D(
        PTstCtrl_C_3), .Y(n1511) );
    zor4b U429 ( .A(TEST_FORCE_ENABLE), .B(SLAVEMODE), .C(n1495), .D(RUN), .Y(
        n1519) );
    znd2b U430 ( .A(DMA_IDLE4), .B(TD_IDLE4), .Y(n1500) );
    znd2b U431 ( .A(DMA_IDLE3), .B(TD_IDLE3), .Y(n1506) );
    znd2b U432 ( .A(TD_IDLE2), .B(DMA_IDLE2), .Y(n1501) );
    znd3b U433 ( .A(DMA_IDLE1), .B(n1520), .C(TD_IDLE1), .Y(n1496) );
    znr3b U434 ( .A(n1513), .B(n1498), .C(n1517), .Y(n1495) );
    znr3b U435 ( .A(n1521), .B(n1513), .C(n1517), .Y(TEST_FORCE_ENABLE) );
    zan2b U436 ( .A(n1521), .B(n1497), .Y(TEST_K) );
    znr3b U437 ( .A(n1521), .B(n1508), .C(n1517), .Y(TEST_J) );
    zivb U438 ( .A(n1498), .Y(n1521) );
    zivb U439 ( .A(n1508), .Y(n1513) );
    zivb U440 ( .A(n1499), .Y(n1520) );
    zind2b U441 ( .A(DBG_GO), .B(DBG_IDLE), .Y(n1502) );
    zivb U442 ( .A(n1510), .Y(n1514) );
    zdffqsb_ DBG_PCLK_EN_2T_reg ( .CK(PCLK66), .D(DBG_PCLK_EN_T), .S(HRST_), 
        .Q(DBG_PCLK_EN_2T) );
    zdffqsb_ DMA_CLK60M_EN1_P_reg ( .CK(CLK60M), .D(DMA_CLK60M_EN1_P1171), .S(
        HRST_), .Q(DMA_CLK60M_EN1_P) );
    zdffqsb_ EHCIFLOW_PCLK_EN_P_reg ( .CK(PCLK66), .D(EHCIFLOW_PCLK_EN_P501), 
        .S(HRST_), .Q(EHCIFLOW_PCLK_EN_P) );
    zdffqsb_ EHCI_DMA_EN4_P_reg ( .CK(PCLK66), .D(EHCI_DMA_EN4_P887), .S(HRST_
        ), .Q(EHCI_DMA_EN4_P) );
    zdffqsb_ EHCI_DMA_EN3_2T_reg ( .CK(PCLK66), .D(EHCI_DMA_EN3_T), .S(HRST_), 
        .Q(EHCI_DMA_EN3_2T) );
    zdffqsb_ HS_MAC_TX_EN_2T_reg ( .CK(CLK60M), .D(HS_MAC_TX_EN_T), .S(HRST_), 
        .Q(HS_MAC_TX_EN_2T) );
    zdffqsb_ EHCI_DMA_EN4_T_reg ( .CK(PCLK66), .D(EHCI_DMA_EN4_P), .S(HRST_), 
        .Q(EHCI_DMA_EN4_T) );
    zdffqsb_ EHCIFLOW_PCLK_EN_2T_reg ( .CK(PCLK66), .D(EHCIFLOW_PCLK_EN_T), 
        .S(HRST_), .Q(EHCIFLOW_PCLK_EN_2T) );
    zdffqsb_ EHCIFLOW_PCLK_EN_T_reg ( .CK(PCLK66), .D(EHCIFLOW_PCLK_EN_P), .S(
        HRST_), .Q(EHCIFLOW_PCLK_EN_T) );
    zdffqsb_ EHCI_DMA_EN2_T_reg ( .CK(PCLK66), .D(EHCI_DMA_EN2_P), .S(HRST_), 
        .Q(EHCI_DMA_EN2_T) );
    zdffqsb_ EHCI_DMA_EN1_2T_reg ( .CK(PCLK66), .D(EHCI_DMA_EN1_T), .S(HRST_), 
        .Q(EHCI_DMA_EN1_2T) );
    zdffqsb_ EHCI_DMA_EN3_T_reg ( .CK(PCLK66), .D(EHCI_DMA_EN3_P), .S(HRST_), 
        .Q(EHCI_DMA_EN3_T) );
    zdffqsb_ EHCI_DMA_EN3_P_reg ( .CK(PCLK66), .D(EHCI_DMA_EN3_P881), .S(HRST_
        ), .Q(EHCI_DMA_EN3_P) );
    zdffqsb_ EHCI_DMA_EN2_P_reg ( .CK(PCLK66), .D(EHCI_DMA_EN2_P875), .S(HRST_
        ), .Q(EHCI_DMA_EN2_P) );
    zdffqsb_ MAC_CLK60M_EN_2T_reg ( .CK(CLK60M), .D(MAC_CLK60M_EN_T), .S(HRST_
        ), .Q(MAC_CLK60M_EN_2T) );
    zdffqsb_ HS_MAC_RX_EN_2T_reg ( .CK(CLK60M), .D(HS_MAC_RX_EN_T), .S(HRST_), 
        .Q(HS_MAC_RX_EN_2T) );
    zdffqsb_ DMA_CLK60M_EN2_P_reg ( .CK(CLK60M), .D(DMA_CLK60M_EN2_P1177), .S(
        HRST_), .Q(DMA_CLK60M_EN2_P) );
    zdffqsb_ EHCI_DMA_EN4_2T_reg ( .CK(PCLK66), .D(EHCI_DMA_EN4_T), .S(HRST_), 
        .Q(EHCI_DMA_EN4_2T) );
    zdffqsb_ DMA_CLK60M_EN3_P_reg ( .CK(CLK60M), .D(DMA_CLK60M_EN3_P1183), .S(
        HRST_), .Q(DMA_CLK60M_EN3_P) );
    zdffqsb_ HS_MAC_TX_EN_P_reg ( .CK(CLK60M), .D(HS_MAC_TX_EN_P701), .S(HRST_
        ), .Q(HS_MAC_TX_EN_P) );
    zdffqsb_ HS_MAC_RX_EN_P_reg ( .CK(CLK60M), .D(HS_MAC_RX_EN_P771), .S(HRST_
        ), .Q(HS_MAC_RX_EN_P) );
    zdffqsb_ DBG_PCLK_EN_P_reg ( .CK(PCLK66), .D(DBG_PCLK_EN_P1321), .S(HRST_), 
        .Q(DBG_PCLK_EN_P) );
    zdffqsb_ MAC_CLK60M_EN_T_reg ( .CK(CLK60M), .D(MAC_CLK60M_EN_P), .S(HRST_), 
        .Q(MAC_CLK60M_EN_T) );
    zdffqsb_ DMA_CLK60M_EN4_P_reg ( .CK(CLK60M), .D(DMA_CLK60M_EN4_P1189), .S(
        HRST_), .Q(DMA_CLK60M_EN4_P) );
    zdffqsb_ EHCI_DMA_EN1_P_reg ( .CK(PCLK66), .D(EHCI_DMA_EN1_P869), .S(HRST_
        ), .Q(EHCI_DMA_EN1_P) );
    zdffqsb_ EHCI_DMA_EN1_T_reg ( .CK(PCLK66), .D(EHCI_DMA_EN1_P), .S(HRST_), 
        .Q(EHCI_DMA_EN1_T) );
    zdffqsb_ MAC_CLK60M_EN_P_reg ( .CK(CLK60M), .D(MAC_CLK60M_EN_P593), .S(
        HRST_), .Q(MAC_CLK60M_EN_P) );
    zdffqsb_ DBG_PCLK_EN_T_reg ( .CK(PCLK66), .D(DBG_PCLK_EN_P), .S(HRST_), 
        .Q(DBG_PCLK_EN_T) );
    zdffqsb_ EHCI_DMA_EN2_2T_reg ( .CK(PCLK66), .D(EHCI_DMA_EN2_T), .S(HRST_), 
        .Q(EHCI_DMA_EN2_2T) );
    zdffqsb_ HS_MAC_RX_EN_T_reg ( .CK(CLK60M), .D(HS_MAC_RX_EN_P), .S(HRST_), 
        .Q(HS_MAC_RX_EN_T) );
    zdffqsb_ HS_MAC_TX_EN_T_reg ( .CK(CLK60M), .D(HS_MAC_TX_EN_P), .S(HRST_), 
        .Q(HS_MAC_TX_EN_T) );
endmodule


module HS_SYNC66 ( PCLK66, HRST_, RUN_C, RUN_C_66, HSERR_S, HSERR_S_66, 
    BIST_RUN_C, BIST_RUN_C_66, BIST_ERR_S, BIST_ERR_S_66, ERRINT_S, 
    ERRINT_S_66, USBINT_S, USBINT_S_66, MABORT, MABORT_66, TABORT, TABORT_66, 
    ROLLOVER_S, ROLLOVER_S_66, INTASYNC_S, INTASYNC_S_66, PORTCHG_S, 
    PORTCHG_S_66, FRNUM_PCLK_LATCH, FRNUM_PCLK_LATCH_66, DBG_COMPL, 
    DBG_COMPL_66, SYNC_SPAREA, SYNC_SPAREA_66, SYNC_SPAREB, SYNC_SPAREB_66 );
input  PCLK66, HRST_, RUN_C, HSERR_S, BIST_RUN_C, BIST_ERR_S, ERRINT_S, 
    USBINT_S, MABORT, TABORT, ROLLOVER_S, INTASYNC_S, PORTCHG_S, 
    FRNUM_PCLK_LATCH, DBG_COMPL, SYNC_SPAREA, SYNC_SPAREB;
output RUN_C_66, HSERR_S_66, BIST_RUN_C_66, BIST_ERR_S_66, ERRINT_S_66, 
    USBINT_S_66, MABORT_66, TABORT_66, ROLLOVER_S_66, INTASYNC_S_66, 
    PORTCHG_S_66, FRNUM_PCLK_LATCH_66, DBG_COMPL_66, SYNC_SPAREA_66, 
    SYNC_SPAREB_66;
    wire SYNC_SPAREA2, MABORT3, SPAREO6, DBG_COMPL3, USBINT_S3, PORTCHG_S2, 
        HSERR_S2, SPAREO0_, ROLLOVER_S2, SPAREO1, HSERR_S3, PORTCHG_S3, 
        SPAREO0, ROLLOVER_S3, DBG_COMPL2, MABORT2, SPAREO7, SYNC_SPAREA3, 
        USBINT_S2, SPAREO5, TABORT2, RUN_C3, SYNC_SPAREB3, ERRINT_S2, 
        BIST_RUN_C2, INTASYNC_S2, SPAREO2, FRNUM_PCLK_LATCH3, BIST_ERR_S2, 
        INTASYNC_S3, BIST_RUN_C3, SYNC_SPAREB2, ERRINT_S3, BIST_ERR_S3, 
        SPAREO3, SPAREO1_, FRNUM_PCLK_LATCH2, RUN_C2, TABORT3, SPAREO4;
    zivb SPARE366 ( .A(SPAREO5), .Y(SPAREO6) );
    zdffrb SPARE361 ( .CK(PCLK66), .D(SPAREO7), .R(1'b1), .Q(SPAREO1), .QN(
        SPAREO1_) );
    zdffrb SPARE360 ( .CK(PCLK66), .D(1'b0), .R(1'b1), .Q(SPAREO0), .QN(
        SPAREO0_) );
    znd3b SPARE367 ( .A(SPAREO3), .B(SPAREO6), .C(1'b1), .Y(SPAREO7) );
    zivb SPARE365 ( .A(SPAREO4), .Y(SPAREO5) );
    zaoi211b SPARE362 ( .A(SPAREO0), .B(PORTCHG_S2), .C(SPAREO1_), .D(1'b0), 
        .Y(SPAREO2) );
    zoai21b SPARE363 ( .A(SPAREO1), .B(INTASYNC_S2), .C(1'b1), .Y(SPAREO3) );
    znr3b SPARE364 ( .A(SPAREO2), .B(RUN_C2), .C(SPAREO0_), .Y(SPAREO4) );
    zdffqrb DBG_COMPL2_reg ( .CK(PCLK66), .D(DBG_COMPL), .R(HRST_), .Q(
        DBG_COMPL2) );
    zdffqrb MABORT2_reg ( .CK(PCLK66), .D(MABORT), .R(HRST_), .Q(MABORT2) );
    zdffqrb INTASYNC_S2_reg ( .CK(PCLK66), .D(INTASYNC_S), .R(HRST_), .Q(
        INTASYNC_S2) );
    zdffqrb_ FRNUM_PCLK_LATCH3_reg ( .CK(PCLK66), .D(FRNUM_PCLK_LATCH2), .R(
        HRST_), .Q(FRNUM_PCLK_LATCH3) );
    zdffqrb_ PORTCHG_S3_reg ( .CK(PCLK66), .D(PORTCHG_S2), .R(HRST_), .Q(
        PORTCHG_S3) );
    zdffqrb_ SYNC_SPAREB3_reg ( .CK(PCLK66), .D(SYNC_SPAREB2), .R(HRST_), .Q(
        SYNC_SPAREB3) );
    zdffqrb_ TABORT3_reg ( .CK(PCLK66), .D(TABORT2), .R(HRST_), .Q(TABORT3) );
    zdffqrb_ BIST_ERR_S3_reg ( .CK(PCLK66), .D(BIST_ERR_S2), .R(HRST_), .Q(
        BIST_ERR_S3) );
    zdffqrb ROLLOVER_S2_reg ( .CK(PCLK66), .D(ROLLOVER_S), .R(HRST_), .Q(
        ROLLOVER_S2) );
    zdffqrb USBINT_S2_reg ( .CK(PCLK66), .D(USBINT_S), .R(HRST_), .Q(USBINT_S2
        ) );
    zdffqrb_ BIST_RUN_C3_reg ( .CK(PCLK66), .D(BIST_RUN_C2), .R(HRST_), .Q(
        BIST_RUN_C3) );
    zdffqrb RUN_C2_reg ( .CK(PCLK66), .D(RUN_C), .R(HRST_), .Q(RUN_C2) );
    zdffqrb SYNC_SPAREA2_reg ( .CK(PCLK66), .D(SYNC_SPAREA), .R(HRST_), .Q(
        SYNC_SPAREA2) );
    zdffqrb_ ERRINT_S3_reg ( .CK(PCLK66), .D(ERRINT_S2), .R(HRST_), .Q(
        ERRINT_S3) );
    zdffqrb HSERR_S2_reg ( .CK(PCLK66), .D(HSERR_S), .R(HRST_), .Q(HSERR_S2)
         );
    zdffqrb BIST_RUN_C2_reg ( .CK(PCLK66), .D(BIST_RUN_C), .R(HRST_), .Q(
        BIST_RUN_C2) );
    zdffqrb_ USBINT_S3_reg ( .CK(PCLK66), .D(USBINT_S2), .R(HRST_), .Q(
        USBINT_S3) );
    zdffqrb_ RUN_C3_reg ( .CK(PCLK66), .D(RUN_C2), .R(HRST_), .Q(RUN_C3) );
    zdffqrb_ SYNC_SPAREA3_reg ( .CK(PCLK66), .D(SYNC_SPAREA2), .R(HRST_), .Q(
        SYNC_SPAREA3) );
    zdffqrb ERRINT_S2_reg ( .CK(PCLK66), .D(ERRINT_S), .R(HRST_), .Q(ERRINT_S2
        ) );
    zdffqrb_ HSERR_S3_reg ( .CK(PCLK66), .D(HSERR_S2), .R(HRST_), .Q(HSERR_S3)
         );
    zdffqrb_ DBG_COMPL3_reg ( .CK(PCLK66), .D(DBG_COMPL2), .R(HRST_), .Q(
        DBG_COMPL3) );
    zdffqrb_ MABORT3_reg ( .CK(PCLK66), .D(MABORT2), .R(HRST_), .Q(MABORT3) );
    zdffqrb_ INTASYNC_S3_reg ( .CK(PCLK66), .D(INTASYNC_S2), .R(HRST_), .Q(
        INTASYNC_S3) );
    zdffqrb PORTCHG_S2_reg ( .CK(PCLK66), .D(PORTCHG_S), .R(HRST_), .Q(
        PORTCHG_S2) );
    zdffqrb FRNUM_PCLK_LATCH2_reg ( .CK(PCLK66), .D(FRNUM_PCLK_LATCH), .R(
        HRST_), .Q(FRNUM_PCLK_LATCH2) );
    zdffqrb SYNC_SPAREB2_reg ( .CK(PCLK66), .D(SYNC_SPAREB), .R(HRST_), .Q(
        SYNC_SPAREB2) );
    zdffqrb TABORT2_reg ( .CK(PCLK66), .D(TABORT), .R(HRST_), .Q(TABORT2) );
    zdffqrb BIST_ERR_S2_reg ( .CK(PCLK66), .D(BIST_ERR_S), .R(HRST_), .Q(
        BIST_ERR_S2) );
    zdffqrb_ ROLLOVER_S3_reg ( .CK(PCLK66), .D(ROLLOVER_S2), .R(HRST_), .Q(
        ROLLOVER_S3) );
    zor3b U186 ( .A(DBG_COMPL3), .B(DBG_COMPL), .C(DBG_COMPL2), .Y(
        DBG_COMPL_66) );
    zor3b U187 ( .A(INTASYNC_S3), .B(INTASYNC_S), .C(INTASYNC_S2), .Y(
        INTASYNC_S_66) );
    zor3b U188 ( .A(BIST_ERR_S3), .B(BIST_ERR_S), .C(BIST_ERR_S2), .Y(
        BIST_ERR_S_66) );
    zor3b U189 ( .A(ROLLOVER_S3), .B(ROLLOVER_S), .C(ROLLOVER_S2), .Y(
        ROLLOVER_S_66) );
    zor3b U190 ( .A(FRNUM_PCLK_LATCH), .B(FRNUM_PCLK_LATCH2), .C(
        FRNUM_PCLK_LATCH3), .Y(FRNUM_PCLK_LATCH_66) );
    zor3b U191 ( .A(ERRINT_S3), .B(ERRINT_S), .C(ERRINT_S2), .Y(ERRINT_S_66)
         );
    zor3b U192 ( .A(USBINT_S), .B(USBINT_S2), .C(USBINT_S3), .Y(USBINT_S_66)
         );
    zor3b U193 ( .A(RUN_C3), .B(RUN_C), .C(RUN_C2), .Y(RUN_C_66) );
    zor3b U194 ( .A(MABORT3), .B(MABORT), .C(MABORT2), .Y(MABORT_66) );
    zor3b U195 ( .A(PORTCHG_S3), .B(PORTCHG_S), .C(PORTCHG_S2), .Y(
        PORTCHG_S_66) );
    zor3b U196 ( .A(HSERR_S3), .B(HSERR_S), .C(HSERR_S2), .Y(HSERR_S_66) );
    zor3b U197 ( .A(SYNC_SPAREB), .B(SYNC_SPAREB2), .C(SYNC_SPAREB3), .Y(
        SYNC_SPAREB_66) );
    zor3b U198 ( .A(TABORT), .B(TABORT2), .C(TABORT3), .Y(TABORT_66) );
    zor3b U199 ( .A(SYNC_SPAREA), .B(SYNC_SPAREA2), .C(SYNC_SPAREA3), .Y(
        SYNC_SPAREA_66) );
    zor3b U200 ( .A(BIST_RUN_C), .B(BIST_RUN_C2), .C(BIST_RUN_C3), .Y(
        BIST_RUN_C_66) );
endmodule


// Verilog netlist generated by Chris Lai, 01/26/2000 (14:06:44)

module HS_USB (UMDATA, ULRDY, UHIT, UFRAMEOE_, UIRDYO_, UADOE_, UFRAMEO_, 
	UIRDYOE_, UCBEOE_, ULOCKOE_, ULOCKO_, /*UPAROE_,*/ TPAROE_,
	UPERROE, UPARO, 
	UPERRO_, UCBE3O_, UCBE2O_, UCBE1O_, UCBE0O_, UINTOE_, UREQO_, USMIO, 
	UAD31O, UAD30O, UAD29O, UAD28O, UAD27O, UAD26O, UAD25O, UAD24O, 
	UAD23O, UAD22O, UAD21O, UAD20O, UAD19O, UAD18O, UAD17O, UAD16O, 
	UAD15O, UAD14O, UAD13O, UAD12O, UAD11O, UAD10O, UAD9O, UAD8O, UAD7O, 
	UAD6O, UAD5O, UAD4O, UAD3O, UAD2O, UAD1O, UAD0O, MA, MWD, MBE_, CREQ,
	MSWR, MRDY_, COMPL, RDYACK,
	/*TESTMIA, MIAT31, 
	MIAT30, MIAT29, MIAT28, MIAT27, MIAT26, MIAT25, MIAT24, MIAT23, 
	MIAT22, MIAT21, MIAT20, MIAT19, MIAT18, MIAT17, MIAT16, MIAT15, 
	MIAT14, MIAT13, MIAT12, MIAT11, MIAT10, MIAT09, MIAT08, MIAT07, 
	MIAT06, MIAT05, MIAT04, MIAT03, MIAT02, MIAT01, MIAT00,*/ UIRQSEL3, 
	UIRQSEL2, UIRQSEL1, UIRQSEL0, /*USBRSM,*/ TRDYI_, IRDYI_, FRAMEI_, 
	STOPI_, DEVSELI_, CBE3I_, CBE2I_, CBE1I_, CBE0I_, AD31I, AD30I, 
	AD29I, AD28I, AD27I, AD26I, AD25I, AD24I, AD23I, AD22I, AD21I, AD20I, 
	AD19I, AD18I, AD17I, AD16I, AD15I, AD14I, AD13I, AD12I, AD11I, AD10I, 
	AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I, SADI, //CLK48, 
	UGNTI_, PCLK, PCLK66, PCLK33_FREE,
	/*PCLK, DP1, DN1, DP2, DN2,*/ UFRMOED_, UCBEOED_, UADOED_, 
	UIRDYED_, UPAROED_, /*OC0I_, OC1I_,*/ PORTDIR1, PORTDIR2, /*RXC1, RXC2, 
	RXD1, RXD2,*/ DEVSELO_, TRDYO_, TRDYOE_, IDSELI, FUNCSEL, PARI, 
	PERRI_, STOPO_, PMSTR, MABORT, TABORT, ENOCPY, OCUPY_SEL, HRST_,
	/*CLK_12MI,*/ HCRESET,
	PORTSC1, PORTSC2, PORTSC3, PORTSC4, PORTSC5, PORTSC6, PORTSC7, PORTSC8,
	CFG_CS, PORTCHG_S,
	PSC_CBE2_A, PSC_CBE1_A, PSC_CBE0_A,
        PSC_CBE2_B, PSC_CBE1_B, PSC_CBE0_B,
        PSC_CBE2_C, PSC_CBE1_C, PSC_CBE0_C,
        PSC_CBE2_D, PSC_CBE1_D, PSC_CBE0_D,
        PSC_CBE2_E, PSC_CBE1_E, PSC_CBE0_E,
        PSC_CBE2_F, PSC_CBE1_F, PSC_CBE0_F,
        PSC_CBE2_G, PSC_CBE1_G, PSC_CBE0_G,
        PSC_CBE2_H, PSC_CBE1_H, PSC_CBE0_H,
	PTstCtrl_A_3, PTstCtrl_A_2, PTstCtrl_A_1, PTstCtrl_A_0,
	PTstCtrl_B_3, PTstCtrl_B_2, PTstCtrl_B_1, PTstCtrl_B_0,
	PTstCtrl_C_3, PTstCtrl_C_2, PTstCtrl_C_1, PTstCtrl_C_0,
	PTstCtrl_D_3, PTstCtrl_D_2, PTstCtrl_D_1, PTstCtrl_D_0,
	PTstCtrl_E_3, PTstCtrl_E_2, PTstCtrl_E_1, PTstCtrl_E_0,
	PTstCtrl_F_3, PTstCtrl_F_2, PTstCtrl_F_1, PTstCtrl_F_0,
	PTstCtrl_G_3, PTstCtrl_G_2, PTstCtrl_G_1, PTstCtrl_G_0,
	PTstCtrl_H_3, PTstCtrl_H_2, PTstCtrl_H_1, PTstCtrl_H_0,
	RxDataOut_A, SquelchOut_A, DisconnectOut_A, TERM_ON_A,
        RxDataOut_B, SquelchOut_B, DisconnectOut_B, TERM_ON_B,
        RxDataOut_C, SquelchOut_C, DisconnectOut_C, TERM_ON_C,
        RxDataOut_D, SquelchOut_D, DisconnectOut_D, TERM_ON_D,
        RxDataOut_E, SquelchOut_E, DisconnectOut_E, TERM_ON_E,
        RxDataOut_F, SquelchOut_F, DisconnectOut_F, TERM_ON_F,
        RxDataOut_G, SquelchOut_G, DisconnectOut_G, TERM_ON_G,
        RxDataOut_H, SquelchOut_H, DisconnectOut_H, TERM_ON_H,
	DIS_TERM_ON_A, DIS_TERM_ON_B, DIS_TERM_ON_C, DIS_TERM_ON_D,
	DIS_TERM_ON_E, DIS_TERM_ON_F, DIS_TERM_ON_G, DIS_TERM_ON_H,
	// USB PME interface
	R61G, R62G, R63G, R84G, R85G,
	FLADJ5, FLADJ4, FLADJ3, FLADJ2, FLADJ1, FLADJ0, ConfigFlag,
	PORTWAKECAP8, PORTWAKECAP7, PORTWAKECAP6, PORTWAKECAP5,
	PORTWAKECAP4, PORTWAKECAP3, PORTWAKECAP2, PORTWAKECAP1, PORTWAKECAP0,
	PWR_STATE1, PWR_STATE0, E_PME_EN, PME_EN, PME_STS, LADO, ADS_PRE,
	PWR_STATE_D0,
	EN_DBG_PORT, DBG_ENABLE_WC, DBG_OWNER, DBG_ENABLE,
	DBG_SEL, DBG_PORT_BLOCKING,
	// USB 2.0 interface
	DATA_TX, TXVALID, TXREADY, RXACTIVE, DATA_RX, TRST_, RXVALID,
	RXSTUFFERR, /*PHYRXERR,*/ RXEOPERR, DIS_STUFF, ASKREPLY, UTM_SOF,
	RCV_POWERUP, TEST_EYE, HS_TRST_,
	// USB PHY option bits
        CP0, CP1, SOF_DISCONN,
        CTRL_A, CTRL_B, CTRL_C, CTRL_D, CTRL_E, CTRL_F, CTRL_G, CTRL_H,
        tst_buferr, loopback, tstmod, rx_block_dis,
        FastLock, LockSpd, TrkSpd, RxDataDly, FastStart, autochk, RDOUT_Enb,
        LBack_Enb, FAST_RST, TMODE, BypassDiv4, UTM_CHKERR,
	sync_fast, sync_jend, SQSET,
	FBABBLE, HCHALT, CLK60M, SetPowner_Dis, PdPHY_Dis, HsEnFB_Dis,
	RVLD, EN_UTM_SPDUP,
	UTM_WR, UTM_DIN, UTM_DOUT,
	/*FOUNDRYID7, FOUNDRYID6, FOUNDRYID5, FOUNDRYID4,
        FOUNDRYID3, FOUNDRYID2, FOUNDRYID1, FOUNDRYID0,*/
	/*EEPHASE, EECFGW0, EECFGW1, EEADO, EECBE, EECS, EESK, EEDI, EEDO,
	EEPA7I, EEPA6I, EEPA5I, EEPA4I, EEPA3I, EEPA2I,*/ EN_EHCI,
	EHCIFLOW_PCLK_EN, MAC_CLK60M_EN, EHCI_DMA_EN1, EHCI_DMA_EN2,
	EHCI_DMA_EN3, EHCI_DMA_EN4, DMA_CLK60M_EN1, DMA_CLK60M_EN2,
	DMA_CLK60M_EN3, DMA_CLK60M_EN4,
	EHCIFLOW_PCLK, MAC_CLK60M, EHCI_DMA1_PCLK, EHCI_DMA2_PCLK,
	EHCI_DMA3_PCLK, EHCI_DMA4_PCLK, DMA1_CLK60M, DMA2_CLK60M,
	DMA3_CLK60M, DMA4_CLK60M,
	EHCIFLOW_CACHE_PCLK, EHCI_DMA1_CACHE_PCLK, EHCI_DMA2_CACHE_PCLK,
	EHCI_DMA3_CACHE_PCLK, EHCI_DMA4_CACHE_PCLK,
	HS_MAC_TX_EN, HS_MAC_RX_EN, HS_MAC_TX_CLK60M, HS_MAC_RX_CLK60M,
	AUTOCHK_CLK60M_EN,
	DBG_PCLK_EN, DBG_CLK60M_EN, DBG_PCLK, DBG_CLK60M,
	CRCERR, PIDERR, TMOUT, TOGMATCH, ENUSB1, ENUSB2, ENUSB3, ENUSB4,
	UMORE, UMORE2LN, TRDYOED_, PCLK33_EN, ATPG_ENI, ATPG_CLK );
input	[7:0]	UTM_WR;
input	[31:0]	UTM_DIN;
output	[63:0]	UTM_DOUT;
output	HS_MAC_TX_EN, HS_MAC_RX_EN, AUTOCHK_CLK60M_EN;
input	HS_MAC_TX_CLK60M, HS_MAC_RX_CLK60M;
output	DBG_PCLK_EN, DBG_CLK60M_EN;
input	DBG_PCLK, DBG_CLK60M;
output	sync_fast, sync_jend;
output	[1:0]	SQSET;
output	EN_UTM_SPDUP;
input	RVLD;
output	EN_DBG_PORT, DBG_ENABLE_WC;
output	DBG_OWNER, DBG_ENABLE, DBG_SEL, DBG_PORT_BLOCKING;
input	PCLK33_FREE;
output	PCLK33_EN;
input	ATPG_CLK;
output	UMORE, UMORE2LN, TRDYOED_;
input	ENUSB1, ENUSB2, ENUSB3, ENUSB4;
output	[31:0]	MA, MWD;
output	[3:0]	MBE_;
output	CREQ, MSWR, MRDY_, COMPL;
input	RDYACK;
input	[31:0]	SADI;
input	EHCIFLOW_PCLK, MAC_CLK60M, EHCI_DMA1_PCLK, EHCI_DMA2_PCLK,
	EHCI_DMA3_PCLK, EHCI_DMA4_PCLK, DMA1_CLK60M, DMA2_CLK60M,
	DMA3_CLK60M, DMA4_CLK60M;
input	EHCIFLOW_CACHE_PCLK, EHCI_DMA1_CACHE_PCLK, EHCI_DMA2_CACHE_PCLK,
	EHCI_DMA3_CACHE_PCLK, EHCI_DMA4_CACHE_PCLK;
output	CRCERR, PIDERR, TMOUT, TOGMATCH;    // output to TEST6~10
output	EHCIFLOW_PCLK_EN, MAC_CLK60M_EN, EHCI_DMA_EN1, EHCI_DMA_EN2,
	EHCI_DMA_EN3, EHCI_DMA_EN4, DMA_CLK60M_EN1, DMA_CLK60M_EN2,
	DMA_CLK60M_EN3, DMA_CLK60M_EN4;
//output	EEPHASE, EECFGW0, EECFGW1, EECS, EESK, EEDI;
input	/*EEDO,*/ EN_EHCI;
//output  [31:0]  EEADO;
//output  [3:0]   EECBE;
//output	EEPA7I, EEPA6I, EEPA5I, EEPA4I, EEPA3I, EEPA2I;
output  CP0, CP1, SOF_DISCONN, loopback, tstmod, rx_block_dis, tst_buferr,
        RDOUT_Enb, FastLock, LBack_Enb, FAST_RST, TMODE, FastStart, BypassDiv4;
output	autochk, SetPowner_Dis, PdPHY_Dis, HsEnFB_Dis;
output  [3:0]   CTRL_A, CTRL_B, CTRL_C, CTRL_D, CTRL_E, CTRL_F, CTRL_G, CTRL_H;
output  [2:0]   RxDataDly;
output  [1:0]   LockSpd, TrkSpd;
output	R61G, R62G, R63G, R84G, R85G, UTM_SOF;
input	FLADJ5, FLADJ4, FLADJ3, FLADJ2, FLADJ1, FLADJ0, ConfigFlag,
	PORTWAKECAP8, PORTWAKECAP7, PORTWAKECAP6, PORTWAKECAP5,
	PORTWAKECAP4, PORTWAKECAP3, PORTWAKECAP2, PORTWAKECAP1, PORTWAKECAP0,
	PWR_STATE1, PWR_STATE0, PME_EN, PME_STS, E_PME_EN, PWR_STATE_D0;
output	ADS_PRE;
output	[31:0]	LADO;
output	[7:0]	DATA_TX;
input	[7:0]	DATA_RX;
output	TRST_, DIS_STUFF, ASKREPLY, RCV_POWERUP, TXVALID;
input	TXREADY, RXACTIVE, RXVALID, RXSTUFFERR, /*PHYRXERR,*/ RXEOPERR, CLK60M;
input	UTM_CHKERR;
input	HS_TRST_;

input	HRST_;//, CLK_12MI;
output	ENOCPY, HCRESET;
output	[1:0] OCUPY_SEL;
output	UMDATA, ULRDY, UHIT, UFRAMEOE_, UIRDYO_, UADOE_, UFRAMEO_, UIRDYOE_;
output	UCBEOE_, ULOCKOE_, ULOCKO_, /*UPAROE_,*/ TPAROE_, UPERROE, UPARO, UPERRO_;
output	UCBE3O_, UCBE2O_, UCBE1O_, UCBE0O_, UINTOE_, UREQO_, USMIO, UAD31O;
output	UAD30O, UAD29O, UAD28O, UAD27O, UAD26O, UAD25O, UAD24O, UAD23O;
output	UAD22O, UAD21O, UAD20O, UAD19O, UAD18O, UAD17O, UAD16O, UAD15O;
output	UAD14O, UAD13O, UAD12O, UAD11O, UAD10O, UAD9O, UAD8O, UAD7O, UAD6O;
output	UAD5O, UAD4O, UAD3O, UAD2O, UAD1O, UAD0O; /*, TESTMIA, MIAT31, MIAT30;
input	MIAT29, MIAT28, MIAT27, MIAT26, MIAT25, MIAT24, MIAT23, MIAT22;
input	MIAT21, MIAT20, MIAT19, MIAT18, MIAT17, MIAT16;
output  MIAT15, MIAT14;
output	MIAT13, MIAT12, MIAT11, MIAT10, MIAT09, MIAT08, MIAT07, MIAT06;
output	MIAT05, MIAT04, MIAT03, MIAT02, MIAT01, MIAT00,*/
output	UIRQSEL3, UIRQSEL2;
output	UIRQSEL1, UIRQSEL0; /*USBRSM,*/ //PMSTR;
input	PMSTR, MABORT, TABORT;
input	TRDYI_, IRDYI_, FRAMEI_, STOPI_, DEVSELI_, CBE3I_, CBE2I_, CBE1I_;
input	CBE0I_, AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I;
input	AD23I, AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, AD14I;
input	AD13I, AD12I, AD11I, AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I;
input	AD2I, AD1I, AD0I, /*CLK48,*/ UGNTI_, PCLK, PCLK66;//PCLK;
//inout	DP1, DN1, DP2, DN2;
output	UFRMOED_, UCBEOED_, UADOED_, UIRDYED_, UPAROED_;
//input	OC0I_, OC1I_;
output	PORTDIR1, PORTDIR2, /*RXC1, RXC2, RXD1, RXD2,*/ DEVSELO_, TRDYO_;
output	TRDYOE_;
input	IDSELI, PARI, PERRI_;
input	[2:0]	FUNCSEL;
output	STOPO_;
input   [31:0]  PORTSC1, PORTSC2, PORTSC3, PORTSC4, PORTSC5, PORTSC6, PORTSC7,
		PORTSC8;
output  CFG_CS;
output	PSC_CBE2_A, PSC_CBE1_A, PSC_CBE0_A,
        PSC_CBE2_B, PSC_CBE1_B, PSC_CBE0_B,
        PSC_CBE2_C, PSC_CBE1_C, PSC_CBE0_C,
        PSC_CBE2_D, PSC_CBE1_D, PSC_CBE0_D,
        PSC_CBE2_E, PSC_CBE1_E, PSC_CBE0_E,
        PSC_CBE2_F, PSC_CBE1_F, PSC_CBE0_F,
        PSC_CBE2_G, PSC_CBE1_G, PSC_CBE0_G,
        PSC_CBE2_H, PSC_CBE1_H, PSC_CBE0_H;
input	PTstCtrl_A_3, PTstCtrl_A_2, PTstCtrl_A_1, PTstCtrl_A_0,
	PTstCtrl_B_3, PTstCtrl_B_2, PTstCtrl_B_1, PTstCtrl_B_0,
	PTstCtrl_C_3, PTstCtrl_C_2, PTstCtrl_C_1, PTstCtrl_C_0,
	PTstCtrl_D_3, PTstCtrl_D_2, PTstCtrl_D_1, PTstCtrl_D_0, PORTCHG_S,
	PTstCtrl_E_3, PTstCtrl_E_2, PTstCtrl_E_1, PTstCtrl_E_0,
	PTstCtrl_F_3, PTstCtrl_F_2, PTstCtrl_F_1, PTstCtrl_F_0,
	PTstCtrl_G_3, PTstCtrl_G_2, PTstCtrl_G_1, PTstCtrl_G_0,
	PTstCtrl_H_3, PTstCtrl_H_2, PTstCtrl_H_1, PTstCtrl_H_0;
output	FBABBLE, HCHALT;
output	DIS_TERM_ON_A, DIS_TERM_ON_B, DIS_TERM_ON_C, DIS_TERM_ON_D,
	DIS_TERM_ON_E, DIS_TERM_ON_F, DIS_TERM_ON_G, DIS_TERM_ON_H;
input	RxDataOut_A, SquelchOut_A, DisconnectOut_A, TERM_ON_A,
        RxDataOut_B, SquelchOut_B, DisconnectOut_B, TERM_ON_B,
        RxDataOut_C, SquelchOut_C, DisconnectOut_C, TERM_ON_C,
        RxDataOut_D, SquelchOut_D, DisconnectOut_D, TERM_ON_D,
        RxDataOut_E, SquelchOut_E, DisconnectOut_E, TERM_ON_E,
        RxDataOut_F, SquelchOut_F, DisconnectOut_F, TERM_ON_F,
        RxDataOut_G, SquelchOut_G, DisconnectOut_G, TERM_ON_G,
        RxDataOut_H, SquelchOut_H, DisconnectOut_H, TERM_ON_H;
output	TEST_EYE;
/*input	FOUNDRYID7, FOUNDRYID6, FOUNDRYID5, FOUNDRYID4,
        FOUNDRYID3, FOUNDRYID2, FOUNDRYID1, FOUNDRYID0;*/
input	ATPG_ENI;	// ATPG enable

wire	[13:0] FRNUM;
//wire	[31:0] PSADO;
wire	[7:0] CACHLN;
wire	[7:0] SOFMOD;
wire	[31:12] FLBASE;
wire	[1:0]   FRLSTSIZE;
wire	[31:0] ASYNCLISTADDR;
wire	[7:0]	INTTHRESHOLD;
wire	[31:0]	SLQUEUEADDR;
wire 	[7:0]	SL_ERROFFSET;
wire	[31:0]	PERIOD_CMD, ASYNC_CMD;
wire	[7:0]	TMOUT_PARM, TXDELAY_PARM;
wire	[3:0]	TURN_PARM;
wire    [31:0]  BIST_PATTERN;
wire    [8:0]   SRAM_ADDR;
wire    [1:0]   SRAM_SEL;
wire    [31:0]  SRAM_RDATA1, SRAM_RDATA2, SRAM_RDATA3, SRAM_RDATA4;
wire [7:0] DBG_BUF_WE;
wire [31:0] DBGPORT_SC, DBGPORT_PID, DBGPORT_ADDR, DBGPORT_BUF1, DBGPORT_BUF2;
wire [7:0] RXPID, DBG_RXPID;
wire [3:0] DBG_RXBCNT;
wire [10:0] RXBCNT;

//wire	[1:0] OCUPY_SEL;

wire VDD = 1'b1;
wire GND = 1'b0;

    /*sivb DNTMIA2 ( .A(VDD), .Y(RSMRSTI) );
    sycbufb TST1 ( .A(MIAT23), .Y(RXC1) );
    sycbufb TST2 ( .A(MIAT22), .Y(RXC2) );
    sycbufb TST3 ( .A(MIAT21), .Y(RXD1) );
    sycbufb TST4 ( .A(MIAT20), .Y(RXD2) );*/
    zivb DNTCLK ( .A(PCLK), .Y(PCICLK_) );
    /*
    USBCLK USBCLK ( .CLKPLL(CLKPLL), .LS(LS), .TRST_(TRST_), .ASKREPLY(
	ASKREPLY), .CLK_12MI(CLK_12MI), .CLK_12M(CLK_12M), .CLK_12M_(CLK_12M_)
	, .CLK_LS(CLK_LS), .CLK_TX_(CLK_TX_), .CLKTXRV(CLKTXRV) );
    */
    zdl1b DNTIRDY ( .A(IRDYI_), .Y(IRDYI_d) );
    zdl1b DNTFRAM ( .A(FRAMEI_), .Y(FRAMEI_d) );

    //san2b DNTCREQ ( .A(CREQ), .B(BMASTREN), .Y(CREQ_GATE) );
    zan2b DNTCREQ ( .A(CREQ_PRE), .B(BMASTREN), .Y(CREQ) );
    zivb DNTUREQ ( .A(CREQ), .Y(UREQO_) );

/*
    UPCIM UPCIM ( .MADDR(MADDR), .MDATA(UMDATA), .UFRAMEOE_(UFRAMEOE_), 
	.UIRDYOE_(UIRDYOE_), .ULOCKOE_(ULOCKOE_), .UCBEOE_(UCBEOE_), .MADOE(
	MADOE), .UPAROE_(UPAROE_), .UPERROE(UPERROE), .UPARO(UPARO), .UPERRO_(
	UPERRO_), .UCBE3O_(UCBE3O_), .UCBE2O_(UCBE2O_), .UCBE1O_(UCBE1O_), 
	.UCBE0O_(UCBE0O_), .UFRAMEO_(UFRAMEO_), .UIRDYO_(UIRDYO_), .UREQO_(
	UREQO_), .ULOCKO_(ULOCKO_), .PMDSEL(PMDSEL), .MABORTS(MABORTS), 
	.TABORTR(TABORTR), .PMSTR(PMSTR), .PERRS(PERRS), .BUSFREE(BUSFREE), 
	.UAD31O(UAD31O), .UAD30O(UAD30O), .UAD29O(UAD29O), .UAD28O(UAD28O), 
	.UAD27O(UAD27O), .UAD26O(UAD26O), .UAD25O(UAD25O), .UAD24O(UAD24O), 
	.UAD23O(UAD23O), .UAD22O(UAD22O), .UAD21O(UAD21O), .UAD20O(UAD20O), 
	.UAD19O(UAD19O), .UAD18O(UAD18O), .UAD17O(UAD17O), .UAD16O(UAD16O), 
	.UAD15O(UAD15O), .UAD14O(UAD14O), .UAD13O(UAD13O), .UAD12O(UAD12O), 
	.UAD11O(UAD11O), .UAD10O(UAD10O), .UAD9O(UAD9O), .UAD8O(UAD8O), 
	.UAD7O(UAD7O), .UAD6O(UAD6O), .UAD5O(UAD5O), .UAD4O(UAD4O), .UAD3O(
	UAD3O), .UAD2O(UAD2O), .UAD1O(UAD1O), .UAD0O(UAD0O), .ADI({AD31I, 
	AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I, AD23I, AD22I, AD21I, 
	AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, AD14I, AD13I, AD12I, AD11I, 
	AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I}), 
	.MSWR(MSWR), .RSTEP(RSTEP), .FB2BKEN(FB2BKEN), .FRAME4(FRAME4), 
	.FRAMEI_(FRAMEI_d), .STOPI_(STOPI_), .LOCKI_(LOCKI_), .TRDYI_(TRDYI_)
	, .IRDYI_(IRDYI_d), .DEVSELI_(DEVSELI_), .CBE3I_(CBE3I_), .CBE2I_(
	CBE2I_), .CBE1I_(CBE1I_), .CBE0I_(CBE0I_), .MBE3_(MBE3_), .MBE2_(MBE2_
	//), .MBE1_(MBE1_), .MBE0_(MBE0_), .CREQ(CREQ), .COMPL(COMPL), .MRDY_(
	), .MBE1_(MBE1_), .MBE0_(MBE0_), .CREQ(CREQ_GATE), .COMPL(COMPL), .MRDY_(
	MRDY_), .CACHEN(CACHEN), .MRDMPLZ(MRDMPLZ), .UGNTI_(UGNTI_), .PCICLK(
	PCLK), .HRST_(HRST_), .UFRMOED_(
	UFRMOED_), .UCBEOED_(UCBEOED_), .UADOED_(UADOED_), .UIRDYED_(UIRDYED_)
	, .UPAROED_(UPAROED_), //.OCUPY_SEL({OCUPY_SEL[1], OCUPY_SEL[0]}), 
	.SERRS(SERRS), .TPAROE_(TPAROE_), .PARI(PARI), .PERRI_(PERRI_), 
	.RPTYERR(RPTYERR), .TDATA(TDATA), .FRAME0(FRAME0), .TGWR(LCMD0), 
	.TRDYO_(TRDYO_), .SERREN(SERREN) );
*/
    HS_SYNC66 HS_SYNC66 ( .PCLK66(PCLK66), .HRST_(HRST_),
        .MABORT(MABORT), .MABORT_66(MABORT_66),
        .TABORT(TABORT), .TABORT_66(TABORT_66),
	.HSERR_S(HSERR_S), .HSERR_S_66(HSERR_S_66),
        .ERRINT_S(ERRINT_S), .ERRINT_S_66(ERRINT_S_66),
        .USBINT_S(USBINT_S), .USBINT_S_66(USBINT_S_66),
	.RUN_C(RUN_C), .RUN_C_66(RUN_C_66),
	.BIST_RUN_C(BIST_RUN_C), .BIST_RUN_C_66(BIST_RUN_C_66),
	.BIST_ERR_S(BIST_ERR_S), .BIST_ERR_S_66(BIST_ERR_S_66),
        .ROLLOVER_S(ROLLOVER_S), .ROLLOVER_S_66(ROLLOVER_S_66),
        .INTASYNC_S(INTASYNC_S), .INTASYNC_S_66(INTASYNC_S_66),
        .PORTCHG_S(PORTCHG_S), .PORTCHG_S_66(PORTCHG_S_66),
	.FRNUM_PCLK_LATCH(FRNUM_PCLK_LATCH),
	.FRNUM_PCLK_LATCH_66(FRNUM_PCLK_LATCH_66),
	.DBG_COMPL(DBG_COMPL), .DBG_COMPL_66(DBG_COMPL_66),
        .SYNC_SPAREA(BIST_ERR_S), .SYNC_SPAREB(USBINT_S) );

    zivb DNTSERR ( .A(VDD), .Y(SERRS) );

    HS_PCIS HS_PCIS ( .PSADO({UAD31O, UAD30O, UAD29O, UAD28O, 
        UAD27O, UAD26O, UAD25O, UAD24O, UAD23O, UAD22O, 
        UAD21O, UAD20O, UAD19O, UAD18O, UAD17O, UAD16O, 
        UAD15O, UAD14O, UAD13O, UAD12O, UAD11O, UAD10O, 
        UAD9O, UAD8O, UAD7O, UAD6O, UAD5O, UAD4O, UAD3O, 
        UAD2O, UAD1O, UAD0O}), .FLBASE({FLBASE[31], FLBASE[30], 
	FLBASE[29], FLBASE[28], FLBASE[27], FLBASE[26], FLBASE[25], FLBASE[24]
	, FLBASE[23], FLBASE[22], FLBASE[21], FLBASE[20], FLBASE[19], 
	FLBASE[18], FLBASE[17], FLBASE[16], FLBASE[15], FLBASE[14], FLBASE[13]
	, FLBASE[12]}), .LIGHTRST(LIGHTRST), .ASYNC_EN(ASYNC_EN),
	.PERIOD_EN(PERIOD_EN), .ASYNC_ACT(ASYNC_ACT), .PERIOD_ACT(PERIOD_ACT),
	.FRLSTSIZE(FRLSTSIZE), .HCRESET(HCRESET), .RUN(RUN),
	.WR_ASYNCADDR(WR_ASYNCADDR), .ASYNCLISTADDR(ASYNCLISTADDR),
	.RECLAMATION(RECLAMATION), .ROLLOVER_S(ROLLOVER_S_66),
	.INTTHRESHOLD(INTTHRESHOLD), /*.IOCSPDINT(IOCSPDINT),
	.USBERRINT(USBERRINT),*/ .ERRINT_EN(ERRINT_EN), .USBINT_EN(USBINT_EN),
	.INTASYNC_EN(INTASYNC_EN), .INTDOORBELL(INTDOORBELL),
	.INTASYNC_S(INTASYNC_S_66), .ASYNCINT(ASYNCINT), .INTASYNC(INTASYNC),
	.SLQUEUEADDR(SLQUEUEADDR), .SLAVEMODE(SLAVEMODE),
	.SLAVE_ACT(SLAVE_ACT), .SL_ERROFFSET(SL_ERROFFSET),
	.CRCERR(CRCERR), .PIDERR(PIDERR), .SL_DATA_PIDERR(SL_DATA_PIDERR),
	.SL_ET_ERR(SL_ET_ERR), .SL_SE_ERR(SL_SE_ERR), .SL_PCIERR(SL_PCIERR),
	.SL_ACK_ERR(SL_ACK_ERR), .SLAVE_ERR(SLAVE_ERR),
	.BIST_RUN(BIST_RUN), .BIST_RUN_C(BIST_RUN_C_66),
        .BIST_ERR_S(BIST_ERR_S_66), .ConfigFlag(ConfigFlag),
	.PORTSC1(PORTSC1), .PORTSC2(PORTSC2), .PORTSC3(PORTSC3),
        .PORTSC4(PORTSC4), .PORTSC5(PORTSC5), .PORTSC6(PORTSC6),
        .PORTSC7(PORTSC7), .PORTSC8(PORTSC8),
	.CFG_CS(CFG_CS), .PORTCHG_S(PORTCHG_S_66),
	.PSC_CBE2_A(PSC_CBE2_A), .PSC_CBE1_A(PSC_CBE1_A),
 	.PSC_CBE0_A(PSC_CBE0_A),
 	.PSC_CBE2_B(PSC_CBE2_B), .PSC_CBE1_B(PSC_CBE1_B),
 	.PSC_CBE0_B(PSC_CBE0_B),
 	.PSC_CBE2_C(PSC_CBE2_C), .PSC_CBE1_C(PSC_CBE1_C),
 	.PSC_CBE0_C(PSC_CBE0_C),
 	.PSC_CBE2_D(PSC_CBE2_D), .PSC_CBE1_D(PSC_CBE1_D),
 	.PSC_CBE0_D(PSC_CBE0_D),
 	.PSC_CBE2_E(PSC_CBE2_E), .PSC_CBE1_E(PSC_CBE1_E),
 	.PSC_CBE0_E(PSC_CBE0_E),
 	.PSC_CBE2_F(PSC_CBE2_F), .PSC_CBE1_F(PSC_CBE1_F),
 	.PSC_CBE0_F(PSC_CBE0_F),
 	.PSC_CBE2_G(PSC_CBE2_G), .PSC_CBE1_G(PSC_CBE1_G),
 	.PSC_CBE0_G(PSC_CBE0_G),
 	.PSC_CBE2_H(PSC_CBE2_H), .PSC_CBE1_H(PSC_CBE1_H),
 	.PSC_CBE0_H(PSC_CBE0_H),

	.R61G(R61G), .R62G(R62G), .R63G(R63G), .R84G(R84G), .R85G(R85G),
	.FLADJ5(FLADJ5), .FLADJ4(FLADJ4), .FLADJ3(FLADJ3), .FLADJ2(FLADJ2),
	.FLADJ1(FLADJ1), .FLADJ0(FLADJ0), .PORTWAKECAP8(PORTWAKECAP8),
	.PORTWAKECAP7(PORTWAKECAP7), .PORTWAKECAP6(PORTWAKECAP6),
	.PORTWAKECAP5(PORTWAKECAP5), .PORTWAKECAP4(PORTWAKECAP4),
	.PORTWAKECAP3(PORTWAKECAP3), .PORTWAKECAP2(PORTWAKECAP2),
	.PORTWAKECAP1(PORTWAKECAP1), .PORTWAKECAP0(PORTWAKECAP0),
	.PWR_STATE1(PWR_STATE1), .PWR_STATE0(PWR_STATE0),
	.PME_EN(PME_EN), .PME_STS(PME_STS), .E_PME_EN(E_PME_EN),
	.PWR_STATE_D0(PWR_STATE_D0),

	.CACHLN({CACHLN[7], CACHLN[6], CACHLN[5], CACHLN[4], 
	CACHLN[3], CACHLN[2], CACHLN[1], CACHLN[0]}), .ULRDY(ULRDY), .UHIT(
	UHIT), .WR_FRNUM(WR_FRNUM), .USBINT(USBINT), .USBEI(USBEI), .USMIO(
	USMIO), .MAXP(MAXP), .SWDBG(SWDBG), .FGR(FGR), .EGSM(EGSM), .GRESET(
	GRESET), .UINTOE_(UINTOE_), .PCI1WAIT(
	PCI1WAIT), .FCFG(FCFG), .PM_EN(PM_EN), .HCISPEC_(HCISPEC_), .PAROPT(
	PAROPT), .BABOPT(BABOPT), .SUSPORT1(SUSPORT1), .PORTRST1(PORTRST1), 
	.RESMPRT1(RESMPRT1), .ENPORT1(ENPORT1), .SUSPORT2(SUSPORT2), 
	.PORTRST2(PORTRST2), .RESMPRT2(RESMPRT2), .ENPORT2(ENPORT2), .FB2BKEN(
	FB2BKEN), .SERREN(SERREN), .RSTEP(RSTEP), .RPTYERR(RPTYERR), .MWRMEN(
	MWRMEN), .CAHCFG_(CAHCFG_), /*.RDYACK(RDYACK),*/ .FRAME0(FRAME0), .FRAME4(
	FRAME4), .SOFMOD({SOFMOD[7], SOFMOD[6], SOFMOD[5], SOFMOD[4], 
	SOFMOD[3], SOFMOD[2], SOFMOD[1], SOFMOD[0]}), .REDUCE(REDUCE), /*.UDIS1(
	UDIS1), .UDIS2(UDIS2), .UENPLL1(UENPLL1), .UENPLL2(UENPLL2), .UPD1(
	UPD1), .UPD2(UPD2), .UTSE01(UTSE01), .UTSE02(UTSE02), .UTXD1(UTXD1), 
	.UTXD2(UTXD2), .UTXE1(UTXE1), .UTXE2(UTXE2), .ULS(ULS), .UCLK48(UCLK48
	), .URST_(URST_), .TESTMIA(TESTMIA),*/ .UIRQSEL3(UIRQSEL3), .UIRQSEL2(
	UIRQSEL2), .UIRQSEL1(UIRQSEL1), .UIRQSEL0(UIRQSEL0), .TESTCNT(TESTCNT)
	, .ENOCPY(ENOCPY), .DISEOP(DISEOP), .DISPRST(DISPRST), .DISSTUFF(
	DISSTUFF), /*.MIAT({MIAT31, MIAT30, MIAT29, MIAT28, MIAT27, MIAT26, 
	MIAT25, MIAT24, MIAT23, MIAT22, MIAT21, MIAT20, MIAT19, MIAT18, MIAT17
	, MIAT16, MIAT15, MIAT14, MIAT13, MIAT12, MIAT11, MIAT10, MIAT09, 
	MIAT08, MIAT07, MIAT06, MIAT05, MIAT04, MIAT03, MIAT02, MIAT01}), */
	/*.ADI({AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I, AD23I, 
	AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, AD14I, AD13I, 
	AD12I, AD11I, AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, 
	//AD1I, AD0I}), .SERRS(SERRS), .PERRS(PERRS), .MABORTS(MABORT), 
	AD1I, AD0I}),*/ .ADI(SADI), .SERRS(SERRS), .PERRS(SERRS),
	.MABORTS(MABORT_66), .TABORTR(TABORT_66),
	.CBE3I_(CBE3I_), .CBE2I_(CBE2I_), .CBE1I_(CBE1I_), 
	.CBE0I_(CBE0I_), .TRDYI_(TRDYI_), .IRDYI_(IRDYI_d), .FRAMEI_(FRAMEI_d)
	, .PMSTR(SERRS), /*.IOCINT(IOCINT), .SPDINT(SPDINT),*/ .ERRINT(ERRINT), 
	/*.FRNUM({FRNUM[15], FRNUM[14], FRNUM[13], FRNUM[12], FRNUM[11], 
	FRNUM[10], FRNUM[9], FRNUM[8], FRNUM[7], FRNUM[6], FRNUM[5], FRNUM[4]
	, FRNUM[3], FRNUM[2], FRNUM[1], FRNUM[0]}),*/ .FRNUM(FRNUM),
	/*.CONN1(MIAT29), .CONN2(MIAT28), .CONNCHG1(CONNCHG1),
	.CONNCHG2(CONNCHG2), .ENCHG1(ENCHG1), 
	.ENCHG2(ENCHG2), .SDP1(MIAT17), .SDP2(MIAT16), .SDN1(MIAT19), .SDN2(
	MIAT18), .LSDEV1(MIAT27), .LSDEV2(MIAT26), .RESMDET1(RESMDET1), 
	.RESMDET2(RESMDET2), .FGREND(FGREND), .SUSACK1(SUSACK1), .RESMEND1(
	RESMEND1), .ENABLE1(ENABLE1), .SUSACK2(SUSACK2), .RESMEND2(RESMEND2), 
	.ENABLE2(ENABLE2), .USBRSM(USBRSM), .OC1I_(OC1I_), .OC0I_(OC0I_),
	.HCHALT_S(HCHALT_S),*/ .HSERR_S(HSERR_S_66), //.PCIERR_S(PCIERR_S), 
	.ERRINT_S(ERRINT_S_66), .USBINT_S(USBINT_S_66), .FATALINT(FATALINT),
	//.RUN_C(RUN_C_66), .CLRHCRST(CLRHCRST), .MAC_EOT(MAC_EOT),
	.RUN_C(RUN_C_66), .CLRHCRST(CLRHCRST), .MAC_EOT(EHCI_DBG_MAC_EOT),
	.PCICLK(PCLK), .HRST_(HRST_),
	.PCICLK_FREE(PCLK33_FREE), .PCIS_ACT(PCIS_ACT),
	/*.CLK_LS(CLK_LS),*/ .OCUPY_SEL({OCUPY_SEL[1], OCUPY_SEL[0]}), 
	.DISTXDLY(DISTXDLY), .DISPFUNDRN(DISPFUNDRN), .ENTXDLY_1(ENTXDLY_1), 
	.ENTXDLY_2(ENTXDLY_2), .ENTXDLY_3(ENTXDLY_3), .SELEOF(SELEOF), 
	.DISTXDLY2(DISTXDLY2), .DISFFCRC0(DISFFCRC0), .DISFFCRC1(DISFFCRC1), 
	.DISPFIFO(DISPFIFO), .DISPFIFO2(DISPFIFO2), .DISRXZERO(DISRXZERO), 
	.ENBMUSMRST(ENBMUSMRST), /*.ENLONGPRESOF(ENLONGPRESOF), .DISFFCRC2(
	DISFFCRC2),*/ .DEVSELI_(DEVSELI_), .DEVSELO_(DEVSELO_), .TRDYO_(TRDYO_)
	, .TRDYOE_(TRDYOE_), .IDSELI(IDSELI), .FUNCSEL(FUNCSEL), .TADOE(TADOE)
	, .TDATA(TDATA), .STOPO_(STOPO_), .TPAROE_(TPAROE_), .LCMD0(LCMD0),
	/*.DISFFCRC3(DISFFCRC3),*/ .DISPSTUFF(DISPSTUFF),
	/*.DISPLATSOF(DISPLATSOF),*/ .DIS_BURST(DIS_BURST),
	.TMOUT_PARM(TMOUT_PARM), .ENISOHANDCHK(ENISOHANDCHK),
	.DISCHKEOPERR(DISCHKEOPERR), .LADO(LADO), .ADS_PRE(ADS_PRE),
	.CP0(CP0), .CP1(CP1), .SOF_DISCONN_CHK(SOF_DISCONN_CHK),
        .CTRL_A(CTRL_A), .CTRL_B(CTRL_B), .CTRL_C(CTRL_C), .CTRL_D(CTRL_D),
	.CTRL_E(CTRL_E), .CTRL_F(CTRL_F), .CTRL_G(CTRL_G), .CTRL_H(CTRL_H),
        .loopback(loopback), .tstmod(tstmod), .rx_block_dis(rx_block_dis),
        .FastLock(FastLock), .LockSpd(LockSpd), .TrkSpd(TrkSpd),
	.sync_fast(sync_fast), .sync_jend(sync_jend), .SQSET(SQSET),
        .RxDataDly(RxDataDly), .RDOUT_Enb(RDOUT_Enb), .LBack_Enb(LBack_Enb),
        .FAST_RST(FAST_RST), .TMODE(TMODE), .BypassDiv4(BypassDiv4),
	.tst_buferr(tst_buferr), .UTM_CHKERR(UTM_CHKERR),
	.TEST_FORCE_ENABLE(TEST_FORCE_ENABLE), .HCHALT(HCHALT),
	.EHCI_IDLE(EHCI_IDLE), .TEST_EYE_EN(TEST_EYE_EN),
	.FastStart(FastStart), .autochk(autochk),
	.RxDataOut_A(RxDataOut_A), .SquelchOut_A(SquelchOut_A),
        .DisconnectOut_A(DisconnectOut_A), .TERM_ON_A(TERM_ON_A),
        .RxDataOut_B(RxDataOut_B), .SquelchOut_B(SquelchOut_B),
        .DisconnectOut_B(DisconnectOut_B), .TERM_ON_B(TERM_ON_B),
        .RxDataOut_C(RxDataOut_C), .SquelchOut_C(SquelchOut_C),
        .DisconnectOut_C(DisconnectOut_C), .TERM_ON_C(TERM_ON_C),
        .RxDataOut_D(RxDataOut_D), .SquelchOut_D(SquelchOut_D),
        .DisconnectOut_D(DisconnectOut_D), .TERM_ON_D(TERM_ON_D),
        .RxDataOut_E(RxDataOut_E), .SquelchOut_E(SquelchOut_E),
        .DisconnectOut_E(DisconnectOut_E), .TERM_ON_E(TERM_ON_E),
        .RxDataOut_F(RxDataOut_F), .SquelchOut_F(SquelchOut_F),
        .DisconnectOut_F(DisconnectOut_F), .TERM_ON_F(TERM_ON_F),
        .RxDataOut_G(RxDataOut_G), .SquelchOut_G(SquelchOut_G),
        .DisconnectOut_G(DisconnectOut_G), .TERM_ON_G(TERM_ON_G),
        .RxDataOut_H(RxDataOut_H), .SquelchOut_H(SquelchOut_H),
        .DisconnectOut_H(DisconnectOut_H), .TERM_ON_H(TERM_ON_H),
	.DIS_TERM_ON_A(DIS_TERM_ON_A), .DIS_TERM_ON_B(DIS_TERM_ON_B),
	.DIS_TERM_ON_C(DIS_TERM_ON_C), .DIS_TERM_ON_D(DIS_TERM_ON_D),
	.DIS_TERM_ON_E(DIS_TERM_ON_E), .DIS_TERM_ON_F(DIS_TERM_ON_F),
	.DIS_TERM_ON_G(DIS_TERM_ON_G), .DIS_TERM_ON_H(DIS_TERM_ON_H),
	.SetPowner_Dis(SetPowner_Dis), .ATPG_ENI(ATPG_ENI),
	.PdPHY_Dis(PdPHY_Dis), .HsEnFB_Dis(HsEnFB_Dis),
	/*.FOUNDRYID0(FOUNDRYID0), .FOUNDRYID1(FOUNDRYID1),
        .FOUNDRYID2(FOUNDRYID2), .FOUNDRYID3(FOUNDRYID3),
        .FOUNDRYID4(FOUNDRYID4), .FOUNDRYID5(FOUNDRYID5),
        .FOUNDRYID6(FOUNDRYID6), .FOUNDRYID7(FOUNDRYID7),*/
	/*.EEPHASE(EEPHASE), .EECFGW0(EECFGW0), .EECFGW1(EECFGW1),
	.EEADO(EEADO), .EECBE(EECBE), .EECS(EECS), .EESK(EESK),
	.EEDI(EEDI), .EEDO(EEDO), .EEPA7I(EEPA7I), .EEPA6I(EEPA6I),
	.EEPA5I(EEPA5I), .EEPA4I(EEPA4I), .EEPA3I(EEPA3I), .EEPA2I(EEPA2I),*/
	.BMASTREN(BMASTREN), .EN_EHCI(EN_EHCI),
	.DISPDRCV(DISPDRCV), .CLKOFF_EN(CLKOFF_EN), .UADS(UADS),
	.TXTMOUT_EN(TXTMOUT_EN),
	.TXDELAY_EN(TXDELAY_EN), .TXDELAY_PARM(TXDELAY_PARM),
	.EN_CHKTOGCRC(EN_CHKTOGCRC), .EN_UTM_RESET(EN_UTM_RESET),
	.TURN_PARM(TURN_PARM), .TRDYOED_(TRDYOED_),
	.ENUSB1(ENUSB1), .ENUSB2(ENUSB2), .ENUSB3(ENUSB3), .ENUSB4(ENUSB4),
	.UTM_RUN(UTM_RUN), .SLEEPTIME_SEL(SLEEPTIME_SEL),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_WR(SRAM_WR), .SRAM_RUN(SRAM_RUN),
        .SRAM_RDATA1(SRAM_RDATA1), .SRAM_RDATA2(SRAM_RDATA2),
        .SRAM_RDATA3(SRAM_RDATA3), .SRAM_RDATA4(SRAM_RDATA4),
	.FRNUM_PCLK_LATCH_66(FRNUM_PCLK_LATCH_66),
	.FORCE_CRCERR(FORCE_CRCERR), .DIS_NARROW_SOF(DIS_NARROW_SOF),
	.DBGPORT_R08G(DBG_BUF_WE[0]), .DBGPORT_R09G(DBG_BUF_WE[1]),
	.DBGPORT_R0AG(DBG_BUF_WE[2]), .DBGPORT_R0BG(DBG_BUF_WE[3]),
        .DBGPORT_R0CG(DBG_BUF_WE[4]), .DBGPORT_R0DG(DBG_BUF_WE[5]),
	.DBGPORT_R0EG(DBG_BUF_WE[6]), .DBGPORT_R0FG(DBG_BUF_WE[7]),
	.EN_DBG_PORT(EN_DBG_PORT), .DBGPORT_SC(DBGPORT_SC),
	.DBGPORT_PID(DBGPORT_PID), .DBGPORT_ADDR(DBGPORT_ADDR),
	.DBGPORT_BUF1(DBGPORT_BUF1), .DBGPORT_BUF2(DBGPORT_BUF2),
        .DBG_COMPL(DBG_COMPL_66), .DBG_XACTERR(DBG_XACTERR),
	.DBG_RXPID(DBG_RXPID), .DBG_RXBCNT(DBG_RXBCNT),
	.DBG_ENABLE_WC(DBG_ENABLE_WC),
	.EN_REF_RVLD(EN_REF_RVLD), .EN_UTM_SPDUP(EN_UTM_SPDUP) );

    zbfd DNT_DBGOWNER ( .A(DBGPORT_SC[30]), .Y(DBG_OWNER) );
    zbfd DNT_DBGENABLE ( .A(DBGPORT_SC[28]), .Y(DBG_ENABLE) );

    //sycbufb DNTMIA ( .A(TESTMIA), .Y(MIAT00) );
    //sycbufb DNTMIA0 ( .A(CLK_12M), .Y(MIAT30) );

//wire BUI_GO2;
//wire #0.5 BUI_GO=BUI_GO2;

    //sdffqa dly6 ( .D(BUI_GO), .CK(PCLK), .Q(BUISTRT) );
    //sycbufb DNTMIA1 ( .A(CLKTXRV), .Y(MIAT31) );
    //sdffqa SYNC01 ( .D(EOT), .CK(PCLK), .Q(EOTQ) );

/*wire HCIADR_31, HCIADR_30, HCIADR_29, HCIADR_28, HCIADR_27, HCIADR_26,
     HCIADR_25, HCIADR_24, HCIADR_23, HCIADR_22, HCIADR_21, HCIADR_20,
     HCIADR_19, HCIADR_18, HCIADR_17, HCIADR_16, HCIADR_15, HCIADR_14,
     HCIADR_13, HCIADR_12, HCIADR_11, HCIADR_10, HCIADR_9, HCIADR_8,
     HCIADR_7, HCIADR_6, HCIADR_5, HCIADR_4, HCIADR_3, HCIADR_2,
     HCIADR_1, HCIADR_0;*/

wire [31:0] HCIADR1, HCIADR2;

/*assign {HCIADR_31, HCIADR_30, HCIADR_29, HCIADR_28, HCIADR_27, HCIADR_26, 
     HCIADR_25, HCIADR_24, HCIADR_23, HCIADR_22, HCIADR_21, HCIADR_20,
     HCIADR_19, HCIADR_18, HCIADR_17, HCIADR_16, HCIADR_15, HCIADR_14,
     HCIADR_13, HCIADR_12, HCIADR_11, HCIADR_10, HCIADR_9, HCIADR_8,
     HCIADR_7, HCIADR_6, HCIADR_5, HCIADR_4, HCIADR_3, HCIADR_2,
     HCIADR_1, HCIADR_0} = HCIADR;*/

/*wire HCIADD_31, HCIADD_30, HCIADD_29, HCIADD_28, HCIADD_27, HCIADD_26,
     HCIADD_25, HCIADD_24, HCIADD_23, HCIADD_22, HCIADD_21, HCIADD_20,
     HCIADD_19, HCIADD_18, HCIADD_17, HCIADD_16, HCIADD_15, HCIADD_14,
     HCIADD_13, HCIADD_12, HCIADD_11, HCIADD_10, HCIADD_9, HCIADD_8,
     HCIADD_7, HCIADD_6, HCIADD_5, HCIADD_4, HCIADD_3, HCIADD_2,
     HCIADD_1, HCIADD_0;*/

wire [31:0] HCIADD1, HCIADD2;

/*assign {HCIADD_31, HCIADD_30, HCIADD_29, HCIADD_28, HCIADD_27, HCIADD_26,
     HCIADD_25, HCIADD_24, HCIADD_23, HCIADD_22, HCIADD_21, HCIADD_20,
     HCIADD_19, HCIADD_18, HCIADD_17, HCIADD_16, HCIADD_15, HCIADD_14,
     HCIADD_13, HCIADD_12, HCIADD_11, HCIADD_10, HCIADD_9, HCIADD_8,
     HCIADD_7, HCIADD_6, HCIADD_5, HCIADD_4, HCIADD_3, HCIADD_2,
     HCIADD_1, HCIADD_0} = HCIADD;*/

//wire BMUSM_RST_EN=0;
//wire DBUFERR=0;
//wire ZEROLEN=0;

wire [10:0] MAXLEN, MAXLEN1, MAXLEN2, MAXLEN3, MAXLEN4, TRAN_MAXLEN1;
wire [31:0] FFRDPCI;
//wire [31:0] BUFPTRA1, BUFPTRA2, BUFPTRB1, BUFPTRB2;
//wire [31:0] BUFPTRC1, BUFPTRC2, BUFPTRD1, BUFPTRD2;
wire [3:0] FBE_;
wire [8:0] FCOUNT;
wire [7:0] HOSTDAT, USBDAT;
wire [7:0] HOSTDAT1, HOSTDAT2, HOSTDAT3, HOSTDAT4, HOSTDAT5;
wire [31:0] WPR1, WPR2, WPR3, WPR4;
wire [7:0] SLADDR;
wire [31:0] MDO, TRAN_BUFPTR1, DMA_BUFPTR1;
wire [19:0] TRAN_BUFPTR2, DMA_BUFPTR2;
//wire SLAVEMODE = 1'b0;

wire [31:0] UADO1, UADO2, UADO3, UADO4;

//assign  UADOE_  = ~(MADOE | TADOE);
    //snr2b DNTUADOE ( .A(MADOE), .B(TADOE), .Y(UADOE_) );
    zivb DNTUADOE ( .A(TADOE), .Y(UADOE_) );

wire [3:0]  PCIDMA_SEL;
wire [4:0]  USBDMA_SEL;
wire [104:0] TRAN_CMD1, TRAN_CMD2, TRAN_CMD3, TRAN_CMD4;
wire [3:0]   ENDP, TXENDP;
wire [6:0]   DEVADDR, TXADDR;
wire [6:0] HUBADDR, HUBPORT;
wire [1:0] SP_ET;
wire [31:0] MA1, MA2, MA3, MA4, MWD1, MWD2, MWD3, MWD4;
wire [51:0] DBG_TRAN_CMD;

    HS_CLKCTL HS_CLKCTL ( .RUN(RUN), .EHCI_IDLE(EHCI_IDLE),
	.USBDMA_SEL(USBDMA_SEL), .SLAVEMODE(SLAVEMODE),
	.TEST_EYE_EN(TEST_EYE_EN), .BIST_RUN(BIST_RUN),
	.HCIREQ1(HCIREQ1), .HCIREQ2(HCIREQ2), .SLHCIREQ(SLHCIREQ),
	.PTstCtrl_A_3(PTstCtrl_A_3), .PTstCtrl_A_2(PTstCtrl_A_2),
        .PTstCtrl_A_1(PTstCtrl_A_1), .PTstCtrl_A_0(PTstCtrl_A_0),
        .PTstCtrl_B_3(PTstCtrl_B_3), .PTstCtrl_B_2(PTstCtrl_B_2),
        .PTstCtrl_B_1(PTstCtrl_B_1), .PTstCtrl_B_0(PTstCtrl_B_0),
        .PTstCtrl_C_3(PTstCtrl_C_3), .PTstCtrl_C_2(PTstCtrl_C_2),
        .PTstCtrl_C_1(PTstCtrl_C_1), .PTstCtrl_C_0(PTstCtrl_C_0),
        .PTstCtrl_D_3(PTstCtrl_D_3), .PTstCtrl_D_2(PTstCtrl_D_2),
        .PTstCtrl_D_1(PTstCtrl_D_1), .PTstCtrl_D_0(PTstCtrl_D_0),
        .PTstCtrl_E_3(PTstCtrl_E_3), .PTstCtrl_E_2(PTstCtrl_E_2),
        .PTstCtrl_E_1(PTstCtrl_E_1), .PTstCtrl_E_0(PTstCtrl_E_0),
        .PTstCtrl_F_3(PTstCtrl_F_3), .PTstCtrl_F_2(PTstCtrl_F_2),
        .PTstCtrl_F_1(PTstCtrl_F_1), .PTstCtrl_F_0(PTstCtrl_F_0),
        .PTstCtrl_G_3(PTstCtrl_G_3), .PTstCtrl_G_2(PTstCtrl_G_2),
        .PTstCtrl_G_1(PTstCtrl_G_1), .PTstCtrl_G_0(PTstCtrl_G_0),
        .PTstCtrl_H_3(PTstCtrl_H_3), .PTstCtrl_H_2(PTstCtrl_H_2),
        .PTstCtrl_H_1(PTstCtrl_H_1), .PTstCtrl_H_0(PTstCtrl_H_0),
	.TD_PARSE_GO1(TD_PARSE_GO1), .TD_PARSE_GO2(TD_PARSE_GO2),
	.TD_PARSE_GO3(TD_PARSE_GO3), .TD_PARSE_GO4(TD_PARSE_GO4),
	.TD_IDLE1(TD_IDLE1), .TD_IDLE2(TD_IDLE2),
	.TD_IDLE3(TD_IDLE3), .TD_IDLE4(TD_IDLE4), .UADS(UADS),
	.EHCIFLOW_PCLK_EN(EHCIFLOW_PCLK_EN),
	.MAC_CLK60M_EN(MAC_CLK60M_EN),
	.EHCI_DMA_EN1(EHCI_DMA_EN1), .EHCI_DMA_EN2(EHCI_DMA_EN2),
	.EHCI_DMA_EN3(EHCI_DMA_EN3), .EHCI_DMA_EN4(EHCI_DMA_EN4),
	.DMA_CLK60M_EN1(DMA_CLK60M_EN1), .DMA_CLK60M_EN2(DMA_CLK60M_EN2),
	.DMA_CLK60M_EN3(DMA_CLK60M_EN3), .DMA_CLK60M_EN4(DMA_CLK60M_EN4),
	.CLKOFF_EN(CLKOFF_EN), .PCLK66(PCLK66), .CLK60M(CLK60M),
	.PCLK33(PCLK33_FREE), .PCIS_ACT(PCIS_ACT), .PCLK33_EN(PCLK33_EN),
	.HRST_(HRST_), .ATPG_ENI(ATPG_ENI),
	.DMA_IDLE1(DMA_IDLE1), .DMA_IDLE2(DMA_IDLE2),
	.DMA_IDLE3(DMA_IDLE3), .DMA_IDLE4(DMA_IDLE4),
	.EN_DBG_PORT(EN_DBG_PORT), .DBG_OWNER(DBG_OWNER),
	.DBG_ENABLE(DBG_ENABLE),
	.DBG_GO(DBGPORT_SC[5]), .DBG_IDLE(DBG_IDLE),
	.DBG_PCLK_EN(DBG_PCLK_EN), .DBG_CLK60M_EN(DBG_CLK60M_EN),
	.TX_PERIOD(TX_PERIOD), .ASKREPLY(ASKREPLY),
	.HS_MAC_TX_EN(HS_MAC_TX_EN), .HS_MAC_RX_EN(HS_MAC_RX_EN),
	.AUTOCHK(autochk), .AUTOCHK_CLK60M_EN(AUTOCHK_CLK60M_EN) );


    HS_DMA_MUX HS_DMA_MUX ( /*.UAD31O(UAD31O), .UAD30O(UAD30O), .UAD29O(UAD29O),
	.UAD28O(UAD28O), .UAD27O(UAD27O), .UAD26O(UAD26O), .UAD25O(UAD25O),
	.UAD24O(UAD24O), .UAD23O(UAD23O), .UAD22O(UAD22O), .UAD21O(UAD21O),
	.UAD20O(UAD20O), .UAD19O(UAD19O), .UAD18O(UAD18O), .UAD17O(UAD17O),
	.UAD16O(UAD16O), .UAD15O(UAD15O), .UAD14O(UAD14O), .UAD13O(UAD13O),
	.UAD12O(UAD12O), .UAD11O(UAD11O), .UAD10O(UAD10O), .UAD9O(UAD9O),
	.UAD8O(UAD8O), .UAD7O(UAD7O), .UAD6O(UAD6O), .UAD5O(UAD5O),
	.UAD4O(UAD4O), .UAD3O(UAD3O), .UAD2O(UAD2O), .UAD1O(UAD1O),
	.UAD0O(UAD0O),
	.UADO1(UADO1), .UADO2(UADO2), .UADO3(UADO3), .UADO4(UADO4),*/
	.MA1(MA1), .MA2(MA2), .MA3(MA3), .MA4(MA4), .MA(MA),
	.MWD1(MWD1), .MWD2(MWD2), .MWD3(MWD3), .MWD4(MWD4), .MWD(MWD),
	.MBE3_(MBE_[3]), .MBE2_(MBE_[2]), .MBE1_(MBE_[1]), .MBE0_(MBE_[0]),
	.MBE3AI_(MBE3AI_), .MBE2AI_(MBE2AI_),
	.MBE1AI_(MBE1AI_), .MBE0AI_(MBE0AI_),
	.MBE3BI_(MBE3BI_), .MBE2BI_(MBE2BI_),
	.MBE1BI_(MBE1BI_), .MBE0BI_(MBE0BI_),
	.MBE3CI_(MBE3CI_), .MBE2CI_(MBE2CI_),
	.MBE1CI_(MBE1CI_), .MBE0CI_(MBE0CI_),
	.MBE3DI_(MBE3DI_), .MBE2DI_(MBE2DI_),
	.MBE1DI_(MBE1DI_), .MBE0DI_(MBE0DI_),
	.CREQ1(CREQ1), .CREQ2(CREQ2), .CREQ3(CREQ3), .CREQ4(CREQ4),
	.CREQ(CREQ_PRE),
	.MRDY1_(MRDY1_), .MRDY2_(MRDY2_), .MRDY3_(MRDY3_), .MRDY4_(MRDY4_),
	.MRDY_(MRDY_),
	.CACHEN1(CACHEN1), .CACHEN2(CACHEN2),
	.CACHEN3(CACHEN3), .CACHEN4(CACHEN4),
	.CACHEN(CACHEN),
	.COMPL1(COMPL1), .COMPL2(COMPL2), .COMPL3(COMPL3), .COMPL4(COMPL4),
	.COMPL(COMPL),
	.MSWR1(MSWR1), .MSWR2(MSWR2), .MSWR3(MSWR3), .MSWR4(MSWR4),
	.MSWR(MSWR),
	.MRDMPLZ1(MRDMPLZ1), .MRDMPLZ2(MRDMPLZ2),
	.MRDMPLZ3(MRDMPLZ3), .MRDMPLZ4(MRDMPLZ4),
	.MRDMPLZ(MRDMPLZ),
	.HOSTDAT1(HOSTDAT1), .HOSTDAT2(HOSTDAT2), .HOSTDAT3(HOSTDAT3),
	.HOSTDAT4(HOSTDAT4), .HOSTDAT5(HOSTDAT5),
	.HOSTDAT(HOSTDAT),
	.LATCHDAT1(LATCHDAT1), .LATCHDAT2(LATCHDAT2),
	.LATCHDAT3(LATCHDAT3), .LATCHDAT4(LATCHDAT4),
	.LATCHDAT5(LATCHDAT5), .LATCHDAT(LATCHDAT),
	.USBPOP1(USBPOP1), .USBPOP2(USBPOP2),
	.USBPOP3(USBPOP3), .USBPOP4(USBPOP4),
	.USBPOP5(USBPOP5), .USBPOP(USBPOP),
	.BUSFREE1(BUSFREE1), .BUSFREE2(BUSFREE2),
	.BUSFREE3(BUSFREE3), .BUSFREE4(BUSFREE4),
	//.BUSFREE(BUSFREE),
	.BUSFREE(1'b1),
	.UGNTI1_(UGNTI1_), .UGNTI2_(UGNTI2_),
	.UGNTI3_(UGNTI3_), .UGNTI4_(UGNTI4_),
	.UGNTI_(UGNTI_),
	.PMDSEL1(PMDSEL1), .PMDSEL2(PMDSEL2),
	.PMDSEL3(PMDSEL3), .PMDSEL4(PMDSEL4),
	//.PMDSEL(PMDSEL),
	.PMDSEL(1'b0),
	.PMSTR1(PMSTR1), .PMSTR2(PMSTR2), .PMSTR3(PMSTR3), .PMSTR4(PMSTR4),
	.PMSTR(PMSTR),
	//.MADDR1(MADDR1), .MADDR2(MADDR2), .MADDR3(MADDR3), .MADDR4(MADDR4),
	//.MADDR(MADDR),
	.MADDR(1'b0),
	.RDYACK1(RDYACK1), .RDYACK2(RDYACK2), .RDYACK3(RDYACK3),
	.RDYACK4(RDYACK4), .RDYACK(RDYACK),
	.MAXLEN(MAXLEN), .TRAN_MAXLEN1(TRAN_MAXLEN1),
	.SLAVE_ACT(SLAVE_ACT), .SLAVEMODE(SLAVEMODE),
	.TEST_PACKET(TEST_PACKET), .SLQUEUEADDR(SLQUEUEADDR),
	.TRAN_BUFPTR1(TRAN_CMD1[103:72]), .TRAN_BUFPTR2(TRAN_CMD1[71:52]),
	.DMA_BUFPTR1(DMA_BUFPTR1), .DMA_BUFPTR2(DMA_BUFPTR2),
	.BIST_ERR_S1(BIST_ERR_S1), .BIST_ERR_S2(BIST_ERR_S2),
	.BIST_ERR_S3(BIST_ERR_S3), .BIST_ERR_S4(BIST_ERR_S4),
	.BIST_ERR_S(BIST_ERR_S),
	//.EOT1(EOT1), .EOT2(EOT2), .EOT3(EOT3), .EOT4(EOT4), .EOT(EOT),
	//.RXERR1(RXERR1), .RXERR2(RXERR2), .RXERR3(RXERR3),
	//.RXERR4(RXERR4), .RXERR(RXERR),
	.TRAN_CMD1(TRAN_CMD1[51:0]), .TRAN_CMD2(TRAN_CMD2[51:0]),
	.TRAN_CMD3(TRAN_CMD3[51:0]), .TRAN_CMD4(TRAN_CMD4[51:0]),
	.TRAN_CMD5(DBG_TRAN_CMD),
	.TXADDR(TXADDR), .TXENDP(TXENDP), .HUBADDR(HUBADDR),
	.HUBPORT(HUBPORT), .SP_SC(SP_SC), .SP_S(SP_S),
	.SP_E(SP_E), .SP_ET(SP_ET), .TD_IN(TD_IN), .TD_OUT(TD_OUT),
	.TD_SETUP(TD_SETUP), .TD_SPLIT(TD_SPLIT), .TD_PING(TD_PING),
	.DAT0(DAT0), .DAT1(DAT1), .DAT2(DAT2), .DATM(DATM),
	.ISO(ISO), .EXEITD(EXEITD),
	.PCIDMA_SEL(PCIDMA_SEL), .USBDMA_SEL(USBDMA_SEL),
	.UMORE1(UMORE1), .UMORE2(UMORE2), .UMORE3(UMORE3), .UMORE4(UMORE4),
	.UMORE2LN1(UMORE2LN1), .UMORE2LN2(UMORE2LN2),
	.UMORE2LN3(UMORE2LN3), .UMORE2LN4(UMORE2LN4),
	.UMORE(UMORE), .UMORE2LN(UMORE2LN),
	.PCICLK(PCLK66), .TRST_(HS_TRST_)
    );

    HS_PER_DMA HS_DMA1 (
	/*.UAD31O(UADO1[31]), .UAD30O(UADO1[30]), .UAD29O(UADO1[29]),
	.UAD28O(UADO1[28]), .UAD27O(UADO1[27]), .UAD26O(UADO1[26]),
	.UAD25O(UADO1[25]), .UAD24O(UADO1[24]), .UAD23O(UADO1[23]),
	.UAD22O(UADO1[22]), .UAD21O(UADO1[21]), .UAD20O(UADO1[20]),
	.UAD19O(UADO1[19]), .UAD18O(UADO1[18]), .UAD17O(UADO1[17]),
	.UAD16O(UADO1[16]), .UAD15O(UADO1[15]), .UAD14O(UADO1[14]),
	.UAD13O(UADO1[13]), .UAD12O(UADO1[12]), .UAD11O(UADO1[11]),
	.UAD10O(UADO1[10]), .UAD9O(UADO1[9]), .UAD8O(UADO1[8]),
	.UAD7O(UADO1[7]), .UAD6O(UADO1[6]), .UAD5O(UADO1[5]),
	.UAD4O(UADO1[4]), .UAD3O(UADO1[3]), .UAD2O(UADO1[2]),
	.UAD1O(UADO1[1]), .UAD0O(UADO1[0]),*/ .MA(MA1), .MWD(MWD1), .WPR(WPR1), 
	.MBE3_(MBE3AI_), .MBE2_(MBE2AI_), .MBE1_(MBE1AI_), .MBE0_(MBE0AI_),
	.CREQ(CREQ1), .MRDY_(MRDY1_), .CACHEN(CACHEN1), .COMPL(COMPL1),
	.MSWR(MSWR1), .MRDMPLZ(MRDMPLZ1), //.XMITNULL(XMITNULL),
	.HCIGNT(HCIGNT1), .TDMAEND(TDMAEND1),
	.TXTHRESH(TXTHRESH1), /*.PSADO31(PSADO[31]), .PSADO30(PSADO[30]), 
	.PSADO29(PSADO[29]), .PSADO28(PSADO[28]), .PSADO27(PSADO[27]), 
	.PSADO26(PSADO[26]), .PSADO25(PSADO[25]), .PSADO24(PSADO[24]), 
	.PSADO23(PSADO[23]), .PSADO22(PSADO[22]), .PSADO21(PSADO[21]), 
	.PSADO20(PSADO[20]), .PSADO19(PSADO[19]), .PSADO18(PSADO[18]), 
	.PSADO17(PSADO[17]), .PSADO16(PSADO[16]), .PSADO15(PSADO[15]), 
	.PSADO14(PSADO[14]), .PSADO13(PSADO[13]), .PSADO12(PSADO[12]), 
	.PSADO11(PSADO[11]), .PSADO10(PSADO[10]), .PSADO9(PSADO[9]),
	.PSADO8(PSADO[8]), .PSADO7(PSADO[7]), .PSADO6(PSADO[6]),
	.PSADO5(PSADO[5]), .PSADO4(PSADO[4]), .PSADO3(PSADO[3]),
	.PSADO2(PSADO[2]), .PSADO1(PSADO[1]), .PSADO0(PSADO[0]),*/
	.AD31I(AD31I), .AD30I(AD30I), .AD29I(AD29I), .AD28I(AD28I),
	.AD27I(AD27I), .AD26I(AD26I), .AD25I(AD25I), .AD24I(AD24I),
	.AD23I(AD23I), .AD22I(AD22I), .AD21I(AD21I), .AD20I(AD20I),
	.AD19I(AD19I), .AD18I(AD18I), .AD17I(AD17I), .AD16I(AD16I),
	.AD15I(AD15I), .AD14I(AD14I), .AD13I(AD13I), .AD12I(AD12I),
	.AD11I(AD11I), .AD10I(AD10I), .AD9I(AD9I), .AD8I(AD8I),
	.AD7I(AD7I), .AD6I(AD6I), .AD5I(AD5I), .AD4I(AD4I),
	.AD3I(AD3I), .AD2I(AD2I), .AD1I(AD1I), .AD0I(AD0I),
	//.BUFPTR1(TRAN_CMD1[115:84]), .BUFPTR2(TRAN_CMD1[83:52]),
	//.BUFPTR1(TRAN_CMD1[103:72]), .BUFPTR2(TRAN_CMD1[71:52]),
	.BUFPTR1(DMA_BUFPTR1), .BUFPTR2(DMA_BUFPTR2),
	//.HCIADR(HCIADR1), .HCIADD(HCIADD1), .MAXLEN(TRAN_CMD1[50:40]),
	.HCIADR(HCIADR1), .HCIADD(HCIADD1), .MAXLEN(TRAN_MAXLEN1),
	.CACHLN7(CACHLN[7]), .CACHLN6(CACHLN[6]), .CACHLN5(CACHLN[5]),
	.CACHLN4(CACHLN[4]), .CACHLN3(CACHLN[3]), .CACHLN2(CACHLN[2]),
	.CACHLN1(CACHLN[1]), .CACHLN0(CACHLN[0]), .CAHCFG_(CAHCFG_),
	.FEMPTY(FEMPTY1), .LATCHDAT(LATCHDAT1), .USBPOP(USBPOP1),
	.USBDAT(USBDAT), .HOSTDAT(HOSTDAT1),
	.QRXERR(RXERR1), .MABORTS(MABORT), .TABORTR(TABORT),
	//.BUSFREE(BUSFREE1), .UGNTI_(UGNTI1_), 
	.BUSFREE(1'b1), .UGNTI_(UGNTI1_), 
	/*.PMDSEL(PMDSEL1),*/ .MWRMEN(MWRMEN), .HCIREQ(HCIREQ1),
	.HCICOMPL(HCICOMPL1), .HCIMWR(HCIMWR1), .HCIMRDY(HCIMRDY1),
	.PMSTR(PMSTR1), .MADDR(MADDR1), .PCI1WAIT(PCI1WAIT), 
	//.EOTQ(EOT1), .IN_DIR(TRAN_CMD1[116]), .RDYACK(RDYACK1), 
	.EOTQ(EOT1), .IN_DIR(TRAN_CMD1[104]), .RDYACK(RDYACK1), 
	/*.UCBE3O_(UCBE3O_), .UCBE2O_(UCBE2O_), .UCBE1O_(UCBE1O_),
	.UCBE0O_(UCBE0O_),*/ .FCFG(FCFG), .HRST_(HRST_),
	.BMUCRST_(BMUCRST_), .DISTXDLY(DISTXDLY), .EOF(EOF),
	.DISTXDLY2(DISTXDLY2), 
	//.BMUSM_RST_EN(BMUSM_RST_EN), .DBUFERR(DBUFERR), .DISPFIFO(DISPFIFO), 
	.BMUSM_RST_EN(1'b0), .DBUFERR(1'b0), .DISPFIFO(DISPFIFO), 
	.DISRXZERO(DISRXZERO), .BUI_GO(BUI_GO1),
	.DISPFIFO2(DISPFIFO2), .ENBMUSMRST(ENBMUSMRST), /*.TADOE(TADOE1),
	.MADOE(MADOE), .UADOE_(UADOE_),*/ //.BOUNDRY(BOUNDRY),
	.TEST_PACKET(TEST_PACKET), .TESTPKTOK(TESTPKTOK),
	.SLAVEMODE(SLAVEMODE), .SLADDR(SLADDR), .DATARDY(DATARDY),
	.SLREAD(SLREAD), .MDO(MDO), .SLAVE_ACT(SLAVE_ACT),
	.BIST_RUN(BIST_RUN), .BIST_RUN_C(BIST_RUN_C),
	.BIST_ERR_S(BIST_ERR_S1), .DIS_BURST(DIS_BURST),
	.PCICLK(EHCI_DMA1_PCLK),
	.HS_TRST_(HS_TRST_), .CLK60M(DMA1_CLK60M), .DMA_IDLE(DMA_IDLE1),
	.UMORE(UMORE1), .UMORE2LN(UMORE2LN1), .ATPG_ENI(ATPG_ENI),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_WR(SRAM_WR), .SRAM_RUN(SRAM_RUN),
        .SRAM_RDATA(SRAM_RDATA1), .SRAM_ID({GND, GND}),
	.ATPG_CLK(ATPG_CLK) );

    HS_PER_DMA HS_DMA2 (
	/*.UAD31O(UADO2[31]), .UAD30O(UADO2[30]), .UAD29O(UADO2[29]),
	.UAD28O(UADO2[28]), .UAD27O(UADO2[27]), .UAD26O(UADO2[26]),
	.UAD25O(UADO2[25]), .UAD24O(UADO2[24]), .UAD23O(UADO2[23]),
	.UAD22O(UADO2[22]), .UAD21O(UADO2[21]), .UAD20O(UADO2[20]),
	.UAD19O(UADO2[19]), .UAD18O(UADO2[18]), .UAD17O(UADO2[17]),
	.UAD16O(UADO2[16]), .UAD15O(UADO2[15]), .UAD14O(UADO2[14]),
	.UAD13O(UADO2[13]), .UAD12O(UADO2[12]), .UAD11O(UADO2[11]),
	.UAD10O(UADO2[10]), .UAD9O(UADO2[9]), .UAD8O(UADO2[8]),
	.UAD7O(UADO2[7]), .UAD6O(UADO2[6]), .UAD5O(UADO2[5]),
	.UAD4O(UADO2[4]), .UAD3O(UADO2[3]), .UAD2O(UADO2[2]),
	.UAD1O(UADO2[1]), .UAD0O(UADO2[0]),*/ .MA(MA2), .MWD(MWD2), .WPR(WPR2), 
	.MBE3_(MBE3BI_), .MBE2_(MBE2BI_), .MBE1_(MBE1BI_), .MBE0_(MBE0BI_),
	.CREQ(CREQ2), .MRDY_(MRDY2_), .CACHEN(CACHEN2), .COMPL(COMPL2),
	.MSWR(MSWR2), .MRDMPLZ(MRDMPLZ2), //.XMITNULL(XMITNULL),
	/*.HCIGNT(HCIGNT),*/ .TDMAEND(TDMAEND2),
	.TXTHRESH(TXTHRESH2), /*.PSADO31(PSADO[31]), .PSADO30(PSADO[30]), 
	.PSADO29(PSADO[29]), .PSADO28(PSADO[28]), .PSADO27(PSADO[27]), 
	.PSADO26(PSADO[26]), .PSADO25(PSADO[25]), .PSADO24(PSADO[24]), 
	.PSADO23(PSADO[23]), .PSADO22(PSADO[22]), .PSADO21(PSADO[21]), 
	.PSADO20(PSADO[20]), .PSADO19(PSADO[19]), .PSADO18(PSADO[18]), 
	.PSADO17(PSADO[17]), .PSADO16(PSADO[16]), .PSADO15(PSADO[15]), 
	.PSADO14(PSADO[14]), .PSADO13(PSADO[13]), .PSADO12(PSADO[12]), 
	.PSADO11(PSADO[11]), .PSADO10(PSADO[10]), .PSADO9(PSADO[9]),
	.PSADO8(PSADO[8]), .PSADO7(PSADO[7]), .PSADO6(PSADO[6]),
	.PSADO5(PSADO[5]), .PSADO4(PSADO[4]), .PSADO3(PSADO[3]),
	.PSADO2(PSADO[2]), .PSADO1(PSADO[1]), .PSADO0(PSADO[0]),*/
	.AD31I(AD31I), .AD30I(AD30I), .AD29I(AD29I), .AD28I(AD28I),
	.AD27I(AD27I), .AD26I(AD26I), .AD25I(AD25I), .AD24I(AD24I),
	.AD23I(AD23I), .AD22I(AD22I), .AD21I(AD21I), .AD20I(AD20I),
	.AD19I(AD19I), .AD18I(AD18I), .AD17I(AD17I), .AD16I(AD16I),
	.AD15I(AD15I), .AD14I(AD14I), .AD13I(AD13I), .AD12I(AD12I),
	.AD11I(AD11I), .AD10I(AD10I), .AD9I(AD9I), .AD8I(AD8I),
	.AD7I(AD7I), .AD6I(AD6I), .AD5I(AD5I), .AD4I(AD4I),
	.AD3I(AD3I), .AD2I(AD2I), .AD1I(AD1I), .AD0I(AD0I),
	//.BUFPTR1(TRAN_CMD2[115:84]), .BUFPTR2(TRAN_CMD2[83:52]),
	.BUFPTR1(TRAN_CMD2[103:72]), .BUFPTR2(TRAN_CMD2[71:52]),
	.HCIADR({32{1'b0}}), .HCIADD({32{1'b0}}), .MAXLEN(TRAN_CMD2[50:40]),
	.CACHLN7(CACHLN[7]), .CACHLN6(CACHLN[6]), .CACHLN5(CACHLN[5]),
	.CACHLN4(CACHLN[4]), .CACHLN3(CACHLN[3]), .CACHLN2(CACHLN[2]),
	.CACHLN1(CACHLN[1]), .CACHLN0(CACHLN[0]), .CAHCFG_(CAHCFG_),
	.FEMPTY(FEMPTY2), .LATCHDAT(LATCHDAT2), .USBPOP(USBPOP2),
	.USBDAT(USBDAT), .HOSTDAT(HOSTDAT2),
	.QRXERR(RXERR2), .MABORTS(MABORT), .TABORTR(TABORT),
	//.BUSFREE(BUSFREE2), .UGNTI_(UGNTI2_), 
	.BUSFREE(1'b1), .UGNTI_(UGNTI2_), 
	/*.PMDSEL(PMDSEL2),*/ .MWRMEN(MWRMEN), .HCIREQ(1'b0), .HCICOMPL(1'b0),
	.HCIMWR(1'b0), .HCIMRDY(1'b0),
	//.PMSTR(PMSTR2), .MADDR(MADDR2), .PCI1WAIT(PCI1WAIT), 
	.PMSTR(PMSTR2), .MADDR(1'b0), .PCI1WAIT(PCI1WAIT), 
	//.EOTQ(EOT2), .IN_DIR(TRAN_CMD2[116]), .RDYACK(RDYACK2), 
	.EOTQ(EOT2), .IN_DIR(TRAN_CMD2[104]), .RDYACK(RDYACK2), 
	/*.UCBE3O_(UCBE3O_), .UCBE2O_(UCBE2O_), .UCBE1O_(UCBE1O_),
	.UCBE0O_(UCBE0O_),*/ .FCFG(FCFG), .HRST_(HRST_),
	.BMUCRST_(BMUCRST_), .DISTXDLY(DISTXDLY), .EOF(EOF),
	.DISTXDLY2(DISTXDLY2), 
	//.BMUSM_RST_EN(BMUSM_RST_EN), .DBUFERR(DBUFERR), .DISPFIFO(DISPFIFO), 
	.BMUSM_RST_EN(1'b0), .DBUFERR(1'b0), .DISPFIFO(DISPFIFO), 
	.DISRXZERO(DISRXZERO), .BUI_GO(BUI_GO2),
	.DISPFIFO2(DISPFIFO2), .ENBMUSMRST(ENBMUSMRST), /*.TADOE(TADOE),
	.MADOE(MADOE), .UADOE_(UADOE_),*/ //.BOUNDRY(BOUNDRY),
	.TEST_PACKET(1'b0), //.TESTPKTOK(TESTPKTOK),
	.SLAVEMODE(1'b0), .SLADDR({8{1'b0}}), //.DATARDY(DATARDY),
	.SLREAD(1'b0), /*.MDO(MDO),*/ .SLAVE_ACT(1'b0),
	.BIST_RUN(BIST_RUN), //.BIST_RUN_C(BIST_RUN_C),
	.BIST_ERR_S(BIST_ERR_S2), .DIS_BURST(DIS_BURST),
	.PCICLK(EHCI_DMA2_PCLK),
	.HS_TRST_(HS_TRST_), .CLK60M(DMA2_CLK60M), .DMA_IDLE(DMA_IDLE2),
	.UMORE(UMORE2), .UMORE2LN(UMORE2LN2), .ATPG_ENI(ATPG_ENI),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_WR(SRAM_WR), .SRAM_RUN(SRAM_RUN),
        .SRAM_RDATA(SRAM_RDATA2), .SRAM_ID({GND, VDD}),
	.ATPG_CLK(ATPG_CLK) );

    HS_ASYNC_DMA HS_DMA3 (
	/*.UAD31O(UADO3[31]), .UAD30O(UADO3[30]), .UAD29O(UADO3[29]),
	.UAD28O(UADO3[28]), .UAD27O(UADO3[27]), .UAD26O(UADO3[26]),
	.UAD25O(UADO3[25]), .UAD24O(UADO3[24]), .UAD23O(UADO3[23]),
	.UAD22O(UADO3[22]), .UAD21O(UADO3[21]), .UAD20O(UADO3[20]),
	.UAD19O(UADO3[19]), .UAD18O(UADO3[18]), .UAD17O(UADO3[17]),
	.UAD16O(UADO3[16]), .UAD15O(UADO3[15]), .UAD14O(UADO3[14]),
	.UAD13O(UADO3[13]), .UAD12O(UADO3[12]), .UAD11O(UADO3[11]),
	.UAD10O(UADO3[10]), .UAD9O(UADO3[9]), .UAD8O(UADO3[8]),
	.UAD7O(UADO3[7]), .UAD6O(UADO3[6]), .UAD5O(UADO3[5]),
	.UAD4O(UADO3[4]), .UAD3O(UADO3[3]), .UAD2O(UADO3[2]),
	.UAD1O(UADO3[1]), .UAD0O(UADO3[0]),*/ .MA(MA3), .MWD(MWD3), .WPR(WPR3), 
	.MBE3_(MBE3CI_), .MBE2_(MBE2CI_), .MBE1_(MBE1CI_), .MBE0_(MBE0CI_),
	.CREQ(CREQ3), .MRDY_(MRDY3_), .CACHEN(CACHEN3), .COMPL(COMPL3),
	.MSWR(MSWR3), .MRDMPLZ(MRDMPLZ3), //.XMITNULL(XMITNULL),
	.HCIGNT(HCIGNT2), .TDMAEND(TDMAEND3),
	.TXTHRESH(TXTHRESH3), /*.PSADO31(PSADO[31]), .PSADO30(PSADO[30]), 
	.PSADO29(PSADO[29]), .PSADO28(PSADO[28]), .PSADO27(PSADO[27]), 
	.PSADO26(PSADO[26]), .PSADO25(PSADO[25]), .PSADO24(PSADO[24]), 
	.PSADO23(PSADO[23]), .PSADO22(PSADO[22]), .PSADO21(PSADO[21]), 
	.PSADO20(PSADO[20]), .PSADO19(PSADO[19]), .PSADO18(PSADO[18]), 
	.PSADO17(PSADO[17]), .PSADO16(PSADO[16]), .PSADO15(PSADO[15]), 
	.PSADO14(PSADO[14]), .PSADO13(PSADO[13]), .PSADO12(PSADO[12]), 
	.PSADO11(PSADO[11]), .PSADO10(PSADO[10]), .PSADO9(PSADO[9]),
	.PSADO8(PSADO[8]), .PSADO7(PSADO[7]), .PSADO6(PSADO[6]),
	.PSADO5(PSADO[5]), .PSADO4(PSADO[4]), .PSADO3(PSADO[3]),
	.PSADO2(PSADO[2]), .PSADO1(PSADO[1]), .PSADO0(PSADO[0]),*/
	.AD31I(AD31I), .AD30I(AD30I), .AD29I(AD29I), .AD28I(AD28I),
	.AD27I(AD27I), .AD26I(AD26I), .AD25I(AD25I), .AD24I(AD24I),
	.AD23I(AD23I), .AD22I(AD22I), .AD21I(AD21I), .AD20I(AD20I),
	.AD19I(AD19I), .AD18I(AD18I), .AD17I(AD17I), .AD16I(AD16I),
	.AD15I(AD15I), .AD14I(AD14I), .AD13I(AD13I), .AD12I(AD12I),
	.AD11I(AD11I), .AD10I(AD10I), .AD9I(AD9I), .AD8I(AD8I),
	.AD7I(AD7I), .AD6I(AD6I), .AD5I(AD5I), .AD4I(AD4I),
	.AD3I(AD3I), .AD2I(AD2I), .AD1I(AD1I), .AD0I(AD0I),
	//.BUFPTR1(TRAN_CMD3[115:84]), .BUFPTR2(TRAN_CMD3[83:52]),
	.BUFPTR1(TRAN_CMD3[103:72]), .BUFPTR2(TRAN_CMD3[71:52]),
	.HCIADR(HCIADR2), .HCIADD(HCIADD2), .MAXLEN(TRAN_CMD3[50:40]),
	.CACHLN7(CACHLN[7]), .CACHLN6(CACHLN[6]), .CACHLN5(CACHLN[5]),
	.CACHLN4(CACHLN[4]), .CACHLN3(CACHLN[3]), .CACHLN2(CACHLN[2]),
	.CACHLN1(CACHLN[1]), .CACHLN0(CACHLN[0]), .CAHCFG_(CAHCFG_),
	.FEMPTY(FEMPTY3), .LATCHDAT(LATCHDAT3), .USBPOP(USBPOP3),
	.USBDAT(USBDAT), .HOSTDAT(HOSTDAT3),
	.QRXERR(RXERR3), .MABORTS(MABORT), .TABORTR(TABORT),
	//.BUSFREE(BUSFREE3), .UGNTI_(UGNTI3_), 
	.BUSFREE(1'b1), .UGNTI_(UGNTI3_), 
	/*.PMDSEL(PMDSEL3),*/ .MWRMEN(MWRMEN), .HCIREQ(HCIREQ2),
	.HCICOMPL(HCICOMPL2), .HCIMWR(HCIMWR2), .HCIMRDY(HCIMRDY2),
	.PMSTR(PMSTR3), .MADDR(MADDR3), .PCI1WAIT(PCI1WAIT), 
	//.EOTQ(EOT3), .IN_DIR(TRAN_CMD3[116]), .RDYACK(RDYACK3), 
	.EOTQ(EOT3), .IN_DIR(TRAN_CMD3[104]), .RDYACK(RDYACK3), 
	/*.UCBE3O_(UCBE3O_), .UCBE2O_(UCBE2O_), .UCBE1O_(UCBE1O_),
	.UCBE0O_(UCBE0O_),*/ .FCFG(FCFG), .HRST_(HRST_),
	.BMUCRST_(BMUCRST_), .DISTXDLY(DISTXDLY), .EOF(EOF),
	.DISTXDLY2(DISTXDLY2), 
	//.BMUSM_RST_EN(BMUSM_RST_EN), .DBUFERR(DBUFERR), .DISPFIFO(DISPFIFO), 
	.BMUSM_RST_EN(1'b0), .DBUFERR(1'b0), .DISPFIFO(DISPFIFO), 
	.DISRXZERO(DISRXZERO), .BUI_GO(BUI_GO3),
	.DISPFIFO2(DISPFIFO2), .ENBMUSMRST(ENBMUSMRST), /*.TADOE(TADOE),
	.MADOE(MADOE), .UADOE_(UADOE_),*/ //.BOUNDRY(BOUNDRY),
	.TEST_PACKET(1'b0), //.TESTPKTOK(TESTPKTOK),
	.SLAVEMODE(1'b0), .SLADDR({8{1'b0}}), //.DATARDY(DATARDY),
	.SLREAD(1'b0), /*.MDO(MDO),*/ .SLAVE_ACT(1'b0),
	.BIST_RUN(BIST_RUN), //.BIST_RUN_C(BIST_RUN_C),
	.BIST_ERR_S(BIST_ERR_S3), .DIS_BURST(DIS_BURST),
	.PCICLK(EHCI_DMA3_PCLK),
	.HS_TRST_(HS_TRST_), .CLK60M(DMA3_CLK60M), .DMA_IDLE(DMA_IDLE3),
	.UMORE(UMORE3), .UMORE2LN(UMORE2LN3), .ATPG_ENI(ATPG_ENI),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_WR(SRAM_WR), .SRAM_RUN(SRAM_RUN),
        .SRAM_RDATA(SRAM_RDATA3), .SRAM_ID({VDD, GND}),
	.ATPG_CLK(ATPG_CLK) );

    HS_ASYNC_DMA HS_DMA4 (
	/*.UAD31O(UADO4[31]), .UAD30O(UADO4[30]), .UAD29O(UADO4[29]),
	.UAD28O(UADO4[28]), .UAD27O(UADO4[27]), .UAD26O(UADO4[26]),
	.UAD25O(UADO4[25]), .UAD24O(UADO4[24]), .UAD23O(UADO4[23]),
	.UAD22O(UADO4[22]), .UAD21O(UADO4[21]), .UAD20O(UADO4[20]),
	.UAD19O(UADO4[19]), .UAD18O(UADO4[18]), .UAD17O(UADO4[17]),
	.UAD16O(UADO4[16]), .UAD15O(UADO4[15]), .UAD14O(UADO4[14]),
	.UAD13O(UADO4[13]), .UAD12O(UADO4[12]), .UAD11O(UADO4[11]),
	.UAD10O(UADO4[10]), .UAD9O(UADO4[9]), .UAD8O(UADO4[8]),
	.UAD7O(UADO4[7]), .UAD6O(UADO4[6]), .UAD5O(UADO4[5]),
	.UAD4O(UADO4[4]), .UAD3O(UADO4[3]), .UAD2O(UADO4[2]),
	.UAD1O(UADO4[1]), .UAD0O(UADO4[0]),*/ .MA(MA4), .MWD(MWD4), .WPR(WPR4), 
	.MBE3_(MBE3DI_), .MBE2_(MBE2DI_), .MBE1_(MBE1DI_), .MBE0_(MBE0DI_),
	.CREQ(CREQ4), .MRDY_(MRDY4_), .CACHEN(CACHEN4), .COMPL(COMPL4),
	.MSWR(MSWR4), .MRDMPLZ(MRDMPLZ4), //.XMITNULL(XMITNULL),
	/*.HCIGNT(HCIGNT),*/ .TDMAEND(TDMAEND4),
	.TXTHRESH(TXTHRESH4), /*.PSADO31(PSADO[31]), .PSADO30(PSADO[30]), 
	.PSADO29(PSADO[29]), .PSADO28(PSADO[28]), .PSADO27(PSADO[27]), 
	.PSADO26(PSADO[26]), .PSADO25(PSADO[25]), .PSADO24(PSADO[24]), 
	.PSADO23(PSADO[23]), .PSADO22(PSADO[22]), .PSADO21(PSADO[21]), 
	.PSADO20(PSADO[20]), .PSADO19(PSADO[19]), .PSADO18(PSADO[18]), 
	.PSADO17(PSADO[17]), .PSADO16(PSADO[16]), .PSADO15(PSADO[15]), 
	.PSADO14(PSADO[14]), .PSADO13(PSADO[13]), .PSADO12(PSADO[12]), 
	.PSADO11(PSADO[11]), .PSADO10(PSADO[10]), .PSADO9(PSADO[9]),
	.PSADO8(PSADO[8]), .PSADO7(PSADO[7]), .PSADO6(PSADO[6]),
	.PSADO5(PSADO[5]), .PSADO4(PSADO[4]), .PSADO3(PSADO[3]),
	.PSADO2(PSADO[2]), .PSADO1(PSADO[1]), .PSADO0(PSADO[0]),*/
	.AD31I(AD31I), .AD30I(AD30I), .AD29I(AD29I), .AD28I(AD28I),
	.AD27I(AD27I), .AD26I(AD26I), .AD25I(AD25I), .AD24I(AD24I),
	.AD23I(AD23I), .AD22I(AD22I), .AD21I(AD21I), .AD20I(AD20I),
	.AD19I(AD19I), .AD18I(AD18I), .AD17I(AD17I), .AD16I(AD16I),
	.AD15I(AD15I), .AD14I(AD14I), .AD13I(AD13I), .AD12I(AD12I),
	.AD11I(AD11I), .AD10I(AD10I), .AD9I(AD9I), .AD8I(AD8I),
	.AD7I(AD7I), .AD6I(AD6I), .AD5I(AD5I), .AD4I(AD4I),
	.AD3I(AD3I), .AD2I(AD2I), .AD1I(AD1I), .AD0I(AD0I),
	//.BUFPTR1(TRAN_CMD4[115:84]), .BUFPTR2(TRAN_CMD4[83:52]),
	.BUFPTR1(TRAN_CMD4[103:72]), .BUFPTR2(TRAN_CMD4[71:52]),
	.HCIADR({32{1'b0}}), .HCIADD({32{1'b0}}), .MAXLEN(TRAN_CMD4[50:40]),
	.CACHLN7(CACHLN[7]), .CACHLN6(CACHLN[6]), .CACHLN5(CACHLN[5]),
	.CACHLN4(CACHLN[4]), .CACHLN3(CACHLN[3]), .CACHLN2(CACHLN[2]),
	.CACHLN1(CACHLN[1]), .CACHLN0(CACHLN[0]), .CAHCFG_(CAHCFG_),
	.FEMPTY(FEMPTY4), .LATCHDAT(LATCHDAT4), .USBPOP(USBPOP4),
	.USBDAT(USBDAT), .HOSTDAT(HOSTDAT4),
	.QRXERR(RXERR4), .MABORTS(MABORT), .TABORTR(TABORT),
	//.BUSFREE(BUSFREE4), .UGNTI_(UGNTI4_), 
	.BUSFREE(1'b1), .UGNTI_(UGNTI4_), 
	/*.PMDSEL(PMDSEL4),*/ .MWRMEN(MWRMEN), .HCIREQ(1'b0), .HCICOMPL(1'b0),
	.HCIMWR(1'b0), .HCIMRDY(1'b0),
	//.PMSTR(PMSTR4), .MADDR(MADDR4), .PCI1WAIT(PCI1WAIT), 
	.PMSTR(PMSTR4), .MADDR(1'b0), .PCI1WAIT(PCI1WAIT), 
	//.EOTQ(EOT4), .IN_DIR(TRAN_CMD4[116]), .RDYACK(RDYACK4), 
	.EOTQ(EOT4), .IN_DIR(TRAN_CMD4[104]), .RDYACK(RDYACK4), 
	/*.UCBE3O_(UCBE3O_), .UCBE2O_(UCBE2O_), .UCBE1O_(UCBE1O_),
	.UCBE0O_(UCBE0O_),*/ .FCFG(FCFG), .HRST_(HRST_),
	.BMUCRST_(BMUCRST_), .DISTXDLY(DISTXDLY), .EOF(EOF),
	.DISTXDLY2(DISTXDLY2), 
	//.BMUSM_RST_EN(BMUSM_RST_EN), .DBUFERR(DBUFERR), .DISPFIFO(DISPFIFO), 
	.BMUSM_RST_EN(1'b0), .DBUFERR(1'b0), .DISPFIFO(DISPFIFO), 
	.DISRXZERO(DISRXZERO), .BUI_GO(BUI_GO4),
	.DISPFIFO2(DISPFIFO2), .ENBMUSMRST(ENBMUSMRST), /*.TADOE(TADOE),
	.MADOE(MADOE), .UADOE_(UADOE_),*/ //.BOUNDRY(BOUNDRY),
	.TEST_PACKET(1'b0), //.TESTPKTOK(TESTPKTOK),
	.SLAVEMODE(1'b0), .SLADDR({8{1'b0}}), //.DATARDY(DATARDY),
	.SLREAD(1'b0), /*.MDO(MDO),*/ .SLAVE_ACT(1'b0),
	.BIST_RUN(BIST_RUN), //.BIST_RUN_C(BIST_RUN_C),
	.BIST_ERR_S(BIST_ERR_S4), .DIS_BURST(DIS_BURST),
	.PCICLK(EHCI_DMA4_PCLK),
	.HS_TRST_(HS_TRST_), .CLK60M(DMA4_CLK60M), .DMA_IDLE(DMA_IDLE4),
	.UMORE(UMORE4), .UMORE2LN(UMORE2LN4), .ATPG_ENI(ATPG_ENI),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_WR(SRAM_WR), .SRAM_RUN(SRAM_RUN),
        .SRAM_RDATA(SRAM_RDATA4), .SRAM_ID({VDD, VDD}),
	.ATPG_CLK(ATPG_CLK) );

    zivb DNTSEL0 ( .A(SELEOF), .Y(SELEOF_) );
    zaoi22b DNTSEL1 ( .A(SELEOF_), .B(EOF1), .C(SELEOF), .D(EOF2), .Y(EOF_) );
    zivb DNTSEL2 ( .A(EOF_), .Y(EOF) );

//wire [5:0]   FLADJ =0;
wire [10:0]  SOFV;
wire [10:0] ACTLEN;

wire [31:0] BUFPTR;

    EHCI EHCI ( .PCI1WAIT(PCI1WAIT), .HCIMRDY1(HCIMRDY1), .HCIMRDY2(HCIMRDY2),
	.RDYACK(RDYACK), .HCICOMPL1(HCICOMPL1), .HCICOMPL2(HCICOMPL2),
        .MABORTS(MABORT), .TABORTR(TABORT),
	.HCIGNT1(HCIGNT1), .HCIGNT2(HCIGNT2), .SLHCIREQ(SLHCIREQ),
	/*.PCICLK(PCLK),*/ .TRST_(HS_TRST_), .PAROPT(PAROPT),
	//.PERRS(PERRS), .SERRS(SERRS), .PMSTR1(PMSTR1), .PMSTR3(PMSTR3),
	.PERRS(SERRS), .SERRS(SERRS), .PMSTR1(PMSTR1), .PMSTR3(PMSTR3),
	.MADDR1(MADDR1), .MADDR3(MADDR3), .UGNTI1_(UGNTI1_), .UGNTI3_(UGNTI3_),
        .ASYNC_EN(ASYNC_EN), .PERIOD_EN(PERIOD_EN),
	.EOF1(EOF1), .EOF2(EOF2), .SOFGEN(SOFGEN),
	.EOFTERM(EOFTERM), .EHCIREQ1(HCIREQ1), .EHCIREQ2(HCIREQ2),
	.FEMPTY1(FEMPTY1), .FEMPTY2(FEMPTY2),
	.FEMPTY3(FEMPTY3), .FEMPTY4(FEMPTY4),
	.ADI({AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I, AD23I,
        AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, AD14I, AD13I,
        AD12I, AD11I, AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I, AD2I,
        AD1I, AD0I}), .SADI(SADI),
	.CLK60M(CLK60M), .FLADJ({FLADJ5, FLADJ4, FLADJ3,
	FLADJ2, FLADJ1, FLADJ0}), .REDUCE(REDUCE),
	.FRNUM(FRNUM), .SOFV(SOFV), .WR_FRNUM(WR_FRNUM),
	.FRLSTSIZE(FRLSTSIZE), .FRNUM_PCLK_LATCH(FRNUM_PCLK_LATCH),
	.RUN(RUN), .HCHALT(HCHALT), .FLBASE(FLBASE),
	.HCIADR1(HCIADR1), .HCIADR2(HCIADR2), .CMDSTART(CMDSTART),
	.MAC_EOT(MAC_EOT),
	.TXSOF(TXSOF), .TDMAEND1(TDMAEND1), .TDMAEND2(TDMAEND2),
	.TDMAEND3(TDMAEND3), .TDMAEND4(TDMAEND4), //.TXTHRESH(TXTHRESH),
	.EOT1(EOT1), .EOT2(EOT2), .EOT3(EOT3), .EOT4(EOT4),
	.CRCERR(CRCERR), .BABBLE(BABBLE), .ACTLEN(ACTLEN),
	.RXERR1(RXERR1), .RXERR2(RXERR2), .RXERR3(RXERR3), .RXERR4(RXERR4),
	.HCIADD1(HCIADD1), .HCIADD2(HCIADD2), .HCIMWR1(HCIMWR1),
	.HCIMWR2(HCIMWR2), .WPR1(WPR1), .WPR2(WPR2), //.BOUNDRY(BOUNDRY),
	.PIDERR(PIDERR), .MAXLEN(MAXLEN),
	.PCIDMA_SEL(PCIDMA_SEL), .USBDMA_SEL(USBDMA_SEL),
	.CREQ1(CREQ1), .CREQ2(CREQ2), .CREQ3(CREQ3), .CREQ4(CREQ4),
	.ASYNCLISTADDR(ASYNCLISTADDR), .TMOUT(TMOUT), .RXNAK(RXNAK),
	.RXNYET(RXNYET), .RXSTALL(RXSTALL), .RXACK(RXACK), .RXDATA0(RXDATA0),
	.RXDATA1(RXDATA1), .RXDATA2(RXDATA2), .RXMDATA(RXMDATA),
	.RXPIDERR(RXPIDERR), .TOGMATCH(TOGMATCH),
	.SPD(SPD),
	.BUI_GO1(BUI_GO1), .BUI_GO2(BUI_GO2), .BUI_GO3(BUI_GO3),
	.BUI_GO4(BUI_GO4),
	.TRAN_CMD1(TRAN_CMD1), .TRAN_CMD2(TRAN_CMD2),
	.TRAN_CMD3(TRAN_CMD3), .TRAN_CMD4(TRAN_CMD4),
	.ASYNC_ACT(ASYNC_ACT), .PERIOD_ACT(PERIOD_ACT), .RUN_C(RUN_C),
	.WR_ASYNCADDR(WR_ASYNCADDR), .RECLAMATION(RECLAMATION),
	.ROLLOVER_S(ROLLOVER_S), .INTTHRESHOLD(INTTHRESHOLD),
	.USBINT(USBINT), .ERRINT(ERRINT), .USBINT_S(USBINT_S),
	.ERRINT_S(ERRINT_S), //.IOCSPDINT(IOCSPDINT), .USBERRINT(USBERRINT),
	.ERRINT_EN(ERRINT_EN), .USBINT_EN(USBINT_EN), .INTASYNC(INTASYNC),
	.INTASYNC_EN(INTASYNC_EN), .INTDOORBELL(INTDOORBELL),
	.INTASYNC_S(INTASYNC_S), .ASYNCINT(ASYNCINT), .EHCIEXE(EHCIEXE),
	.TESTPKTOK(TESTPKTOK), .TEST_PACKET(TEST_PACKET), .SWDBG(SWDBG),
	.HSERR_S(HSERR_S), .SLAVEMODE(SLAVEMODE), //.SLQUEUEADDR(SLQUEUEADDR),
	.SLAVE_ACT(SLAVE_ACT), .BMUCRST_(BMUCRST_), .SLADDR(SLADDR),
	.SLREAD(SLREAD), .DATARDY(DATARDY), .MDO(MDO),
	.PERIOD_CMD(PERIOD_CMD), .ASYNC_CMD(ASYNC_CMD),
	.SL_PERIOD(SL_PERIOD), .SL_DATA_PIDERR(SL_DATA_PIDERR),
	.SL_ET_ERR(SL_ET_ERR), .SL_SE_ERR(SL_SE_ERR),
	.SL_PCIERR(SL_PCIERR), .SL_ACK_ERR(SL_ACK_ERR), .SLAVE_ERR(SLAVE_ERR),
	.SL_ERROFFSET(SL_ERROFFSET), .RXPID(RXPID), .EHCI_IDLE(EHCI_IDLE),
	.TD_IDLE1(TD_IDLE1), .TD_IDLE2(TD_IDLE2),
	.TD_IDLE3(TD_IDLE3), .TD_IDLE4(TD_IDLE4),
	.TD_PARSE_GO1(TD_PARSE_GO1), .TD_PARSE_GO2(TD_PARSE_GO2),
	.TD_PARSE_GO3(TD_PARSE_GO3), .TD_PARSE_GO4(TD_PARSE_GO4),
	.EN_DBG_PORT(EN_DBG_PORT), .DBGPORT_SC(DBGPORT_SC),
	.DBGPORT_PID(DBGPORT_PID), .DBGPORT_ADDR(DBGPORT_ADDR),
        .DBG_COMPL(DBG_COMPL), .DBG_XACTERR(DBG_XACTERR),
	.DBG_RXPID(DBG_RXPID), .DBG_RXBCNT(DBG_RXBCNT),
	.DBG_TRAN_CMD(DBG_TRAN_CMD), .RXBCNT(RXBCNT),
	.EHCIFLOW_PCLK(EHCIFLOW_PCLK), .EHCI_DMA1_PCLK(EHCI_DMA1_PCLK),
	.EHCI_DMA2_PCLK(EHCI_DMA2_PCLK), .EHCI_DMA3_PCLK(EHCI_DMA3_PCLK),
	.EHCI_DMA4_PCLK(EHCI_DMA4_PCLK),
	.EHCIFLOW_CACHE_PCLK(EHCIFLOW_CACHE_PCLK),
	.EHCI_DMA1_CACHE_PCLK(EHCI_DMA1_CACHE_PCLK),
	.EHCI_DMA2_CACHE_PCLK(EHCI_DMA2_CACHE_PCLK),
	.EHCI_DMA3_CACHE_PCLK(EHCI_DMA3_CACHE_PCLK),
	.EHCI_DMA4_CACHE_PCLK(EHCI_DMA4_CACHE_PCLK),
	.SLEEPTIME_SEL(SLEEPTIME_SEL), .DBG_SEL(DBG_SEL),
	.EHCI_DBG_MAC_EOT(EHCI_DBG_MAC_EOT), .DBG_IDLE(DBG_IDLE),
	.DBG_PCLK(DBG_PCLK), .ATPG_ENI(ATPG_ENI) );

//sycbufd DNTBMUCRST ( .A(BMUCRST_), .Y(BMUCRESET_) );

wire [7:0] DATA_TX, DATA_RX;
//wire TEST_J=1'b0;
//wire TEST_K=1'b0;
//assign TEST_PACKET=1'b0;

    HS_MAC HS_MAC ( .DATA_TX(DATA_TX), .TXVALID(TXVALID), .TXREADY(TXREADY),
        .CLK60M(MAC_CLK60M), .TRST_(TRST_), .DIS_STUFF(DIS_STUFF),
        .MAXLEN(MAXLEN), .HOSTDAT(HOSTDAT), .USBPOP(USBPOP),
        .DATA_RX(DATA_RX), .RXACTIVE(RXACTIVE), .RXVALID(RXVALID),
        .USBDAT(USBDAT), .RXEOPERR(RXEOPERR), .RXSTUFFERR(RXSTUFFERR),
        /*.PHYRXERR(PHYRXERR),*/ .DISCHKEOPERR(DISCHKEOPERR),
        .PHYERR(PHYERR), .LATCHDAT(LATCHDAT), //.SLAVEMODE(SLAVEMODE),
        //.TXADDR(DEVADDR), .TXENDP(ENDP), //.FRNUM(FRNUM[10:0]),
        .TXADDR(TXADDR), .TXENDP(TXENDP), //.FRNUM(FRNUM[10:0]),
	.SOFV(SOFV), .HUBADDR(HUBADDR), .EOFTERM(EOFTERM),
        .HUBPORT(HUBPORT), .SP_SC(SP_SC), .SP_S(SP_S), .SP_E(SP_E),
        .SP_ET(SP_ET), .EOF1(EOF1), .EOF2(EOF2), .TD_IN(TD_IN),
        .TD_OUT(TD_OUT), .TD_SETUP(TD_SETUP), .TD_SPLIT(TD_SPLIT),
        .CMDSTART(CMDSTART), .SOFGEN(SOFGEN), .ISO(ISO),
        .DAT0(DAT0), .DAT1(DAT1), .DAT2(DAT2), .DATM(DATM),
        .TMOUT_PARM(TMOUT_PARM), .ASKREPLY(ASKREPLY), .BABBLE(BABBLE),
	.MAC_EOT(MAC_EOT), .TXSOF(TXSOF), .HRST_(HRST_), .HCRESET(HCRESET),
	.CRCERR(CRCERR), .ACTLEN(ACTLEN), .PIDERR(PIDERR), .TMOUT(TMOUT),
	.RXNAK(RXNAK), .RXNYET(RXNYET), .RXSTALL(RXSTALL), .RXACK(RXACK),
	.RXDATA0(RXDATA0), .RXDATA1(RXDATA1), .RXDATA2(RXDATA2),
	.RXMDATA(RXMDATA), .RXPID(RXPID),
	.RXPIDERR(RXPIDERR), .TD_PING(TD_PING), .TOGMATCH(TOGMATCH), .SPD(SPD),
	.LIGHTRST(LIGHTRST), .ENISOHANDCHK(ENISOHANDCHK), .EHCIEXE(1'b0),
	.TEST_J(TEST_J), .TEST_K(TEST_K), .TEST_PACKET(TEST_PACKET),
	.TEST_EYE_EN(TEST_EYE_EN), .TEST_EYE(TEST_EYE),
	.SLAVE_ACT(SLAVE_ACT), .PERIOD_CMD(PERIOD_CMD), .ASYNC_CMD(ASYNC_CMD),
        .SL_PERIOD(SL_PERIOD), .SL_DATA_PIDERR(SL_DATA_PIDERR),
	.SL_ET_ERR(SL_ET_ERR), .SL_SE_ERR(SL_SE_ERR),
	.SL_ACK_ERR(SL_ACK_ERR), .EXEITD(EXEITD),
	.SOF_DISCONN_CHK(SOF_DISCONN_CHK), .SOF_DISCONN(SOF_DISCONN),
	.PTstCtrl_A_3(PTstCtrl_A_3), .PTstCtrl_A_2(PTstCtrl_A_2),
        .PTstCtrl_A_1(PTstCtrl_A_1), .PTstCtrl_A_0(PTstCtrl_A_0),
        .PTstCtrl_B_3(PTstCtrl_B_3), .PTstCtrl_B_2(PTstCtrl_B_2),
        .PTstCtrl_B_1(PTstCtrl_B_1), .PTstCtrl_B_0(PTstCtrl_B_0),
        .PTstCtrl_C_3(PTstCtrl_C_3), .PTstCtrl_C_2(PTstCtrl_C_2),
        .PTstCtrl_C_1(PTstCtrl_C_1), .PTstCtrl_C_0(PTstCtrl_C_0),
        .PTstCtrl_D_3(PTstCtrl_D_3), .PTstCtrl_D_2(PTstCtrl_D_2),
        .PTstCtrl_D_1(PTstCtrl_D_1), .PTstCtrl_D_0(PTstCtrl_D_0),
        .PTstCtrl_E_3(PTstCtrl_E_3), .PTstCtrl_E_2(PTstCtrl_E_2),
        .PTstCtrl_E_1(PTstCtrl_E_1), .PTstCtrl_E_0(PTstCtrl_E_0),
        .PTstCtrl_F_3(PTstCtrl_F_3), .PTstCtrl_F_2(PTstCtrl_F_2),
        .PTstCtrl_F_1(PTstCtrl_F_1), .PTstCtrl_F_0(PTstCtrl_F_0),
        .PTstCtrl_G_3(PTstCtrl_G_3), .PTstCtrl_G_2(PTstCtrl_G_2),
        .PTstCtrl_G_1(PTstCtrl_G_1), .PTstCtrl_G_0(PTstCtrl_G_0),
        .PTstCtrl_H_3(PTstCtrl_H_3), .PTstCtrl_H_2(PTstCtrl_H_2),
        .PTstCtrl_H_1(PTstCtrl_H_1), .PTstCtrl_H_0(PTstCtrl_H_0),
	.TEST_FORCE_ENABLE(TEST_FORCE_ENABLE), .UTM_SOF(UTM_SOF),
	.BABOPT(BABOPT), .FBABBLE(FBABBLE),
	.DISPDRCV(DISPDRCV), .RCV_POWERUP(RCV_POWERUP),
	.TXTMOUT_EN(TXTMOUT_EN),
	.TXDELAY_EN(TXDELAY_EN), .TXDELAY_PARM(TXDELAY_PARM),
	.TURN_PARM(TURN_PARM),
	.ATPG_ENI(ATPG_ENI), .HS_TRST_(HS_TRST_),
	.UTM_RUN(UTM_RUN), .FORCE_CRCERR(FORCE_CRCERR),
	.DIS_NARROW_SOF(DIS_NARROW_SOF), .RXBCNT(RXBCNT),
	.EN_CHKTOGCRC(EN_CHKTOGCRC), .EN_UTM_RESET(EN_UTM_RESET),
	.DBG_TOKEN(DBGPORT_PID[7:0]), .DBG_SENDPID(DBGPORT_PID[15:8]),
	.DBG_SEL(DBG_SEL), .EN_DBG_PORT(EN_DBG_PORT),
	.DBG_PORT_BLOCKING(DBG_PORT_BLOCKING),
	.EN_REF_RVLD(EN_REF_RVLD), .RVLD(RVLD),
	.EN_UTM_SPDUP(EN_UTM_SPDUP), .TX_PERIOD(TX_PERIOD),
	.HS_MAC_TX_CLK60M(HS_MAC_TX_CLK60M),
	.HS_MAC_RX_CLK60M(HS_MAC_RX_CLK60M) );

    DBG_FIFO DBG_FIFO ( .DBG_BUF_WE(DBG_BUF_WE), .DI(LADO),
	.DBGPORT_BUF1(DBGPORT_BUF1), .DBGPORT_BUF2(DBGPORT_BUF2),
	.DBG_GO(DBGPORT_SC[5]), .LATCHDAT(LATCHDAT5),
	.USBPOP(USBPOP5), .USBDAT(USBDAT), .HOSTDAT(HOSTDAT5),
	.UTM_WR(UTM_WR), .UTM_DIN(UTM_DIN), .UTM_DOUT(UTM_DOUT),
	.AUTOCHK(autochk),
	.CLK60M(DBG_CLK60M), .HRST_(HS_TRST_) );

    zivb DNTLOCK ( .A(GND), .Y(LOCKI_) );
    zivb DNTRESP ( .A(VDD), .Y(TRESP) );
    //sdffqa SYNC02 ( .D(RXERR), .CK(PCLK), .Q(QRXERR) );
/*
    MIAMUX MIAMUX ( ._MIARST(MIAT01), .MDIS1(MIAT15), .MDIS2(MIAT14), 
	.MENPLL1(MIAT13), .MENPLL2(MIAT12), .MLS(MIAT03), .MPD1(MIAT11), 
	.MPD2(MIAT10), .MTSE01(MIAT09), .MTSE02(MIAT08), .MTXD1(MIAT07), 
	.MTXD2(MIAT06), .MTXE1(MIAT05), .MTXE2(MIAT04), .MCLK48(MIAT02), 
	.TESTMIA(MIAT00), .TRST_(TRST_), .DIS1(DIS1), .DIS2(DIS2), .ENPLL1(
	ENPLL1), .ENPLL2(ENPLL2), .LS(LS), .PD1(PD1), .PD2(PD2), .TSE01(TSE01)
	, .TSE02(TSE02), .TXD1(TXD1), .TXD2(TXD2), .TXE1(TXE1), .TXE2(TXE2), 
	.CLK48(CLK48), .URST_(URST_), .UDIS1(UDIS1), .UDIS2(UDIS2), .UENPLL1(
	UENPLL1), .UENPLL2(UENPLL2), .ULS(ULS), .UPD1(UPD1), .UPD2(UPD2), 
	.UTSE01(UTSE01), .UTSE02(UTSE02), .UTXD1(UTXD1), .UTXD2(UTXD2), 
	.UTXE1(UTXE1), .UTXE2(UTXE2), .UCLK48(UCLK48) );
*/
    ziva SYNC03 ( .A(VDD), .Y(QRSTPTR) );
    u_redun usb_redun ( .RESET_(HRST_), .CLK(PCLK66), .IN0(AD0I), .IN1(AD1I), 
	.IN2(AD2I), .IN3(AD3I), .IN4(AD4I), .IN5(AD5I), .IN6(AD6I) );
endmodule
 
// USB 2.0 HS periodic DMA controller
module HS_PER_DMA ( /*UAD31O, UAD30O, UAD29O, UAD28O, UAD27O, UAD26O,
		UAD25O, UAD24O, UAD23O, UAD22O, UAD21O, UAD20O,
                UAD19O, UAD18O, UAD17O, UAD16O, UAD15O, UAD14O,
                UAD13O, UAD12O, UAD11O, UAD10O, UAD9O,  UAD8O,
                UAD7O,  UAD6O,  UAD5O,  UAD4O,  UAD3O,  UAD2O,
                UAD1O,  UAD0O,*/
		MA, MWD, WPR,
		MBE3_, MBE2_, MBE1_,MBE0_, CREQ, MRDY_, CACHEN,
		COMPL, MSWR, MRDMPLZ, XMITNULL,
		UMORE, UMORE2LN,
                HCIGNT, TDMAEND, TXTHRESH,
		/*PSADO31, PSADO30, PSADO29, PSADO28, PSADO27, PSADO26,
                PSADO25, PSADO24, PSADO23, PSADO22, PSADO21, PSADO20,
                PSADO19, PSADO18, PSADO17, PSADO16, PSADO15, PSADO14,
                PSADO13, PSADO12, PSADO11, PSADO10, PSADO9,  PSADO8,
                PSADO7,  PSADO6,  PSADO5,  PSADO4,  PSADO3,  PSADO2,
                PSADO1,  PSADO0,*/
		AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I,
		AD23I, AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I,
		AD15I, AD14I, AD13I, AD12I, AD11I, AD10I, AD9I, AD8I,
		AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I,
		BUFPTR1, BUFPTR2, HCIADR, HCIADD, MAXLEN,
		USBDAT, LATCHDAT, USBPOP, HOSTDAT,
		CACHLN7,  CACHLN6,  CACHLN5,  CACHLN4,  CACHLN3,  CACHLN2,
                CACHLN1,  CACHLN0, CAHCFG_,
		FEMPTY,
		QRXERR, MABORTS, TABORTR,
		BUSFREE , UGNTI_, /*PMDSEL,*/ MWRMEN,
		HCIREQ, HCICOMPL, HCIMWR, PMSTR, MADDR, PCI1WAIT,
		EOTQ, IN_DIR, RDYACK,
		//UCBE3O_, UCBE2O_, UCBE1O_,UCBE0O_,
		FCFG, HCIMRDY,
		DISTXDLY, EOF,
		DISTXDLY2, BMUSM_RST_EN, DBUFERR, DISPFIFO,
		DISRXZERO, BUI_GO, DISPFIFO2,
		ENBMUSMRST, /*TADOE, MADOE, UADOE_,*/ BOUNDRY, DIS_BURST,
		TEST_PACKET, SLAVEMODE, SLAVE_ACT, SLADDR, SLREAD,
		BIST_RUN, BIST_RUN_C, BIST_ERR_S, TESTPKTOK, DATARDY,
		MDO, PCICLK, HRST_, BMUCRST_, CLK60M, HS_TRST_, DMA_IDLE,
		ATPG_ENI, BIST_PATTERN, SRAM_ADDR, SRAM_SEL, SRAM_WR, SRAM_RUN,
                SRAM_ID, SRAM_RDATA, ATPG_CLK
		);
input	ATPG_CLK;
input   [31:0]  BIST_PATTERN;
input   [8:0]   SRAM_ADDR;
input   [1:0]   SRAM_SEL, SRAM_ID;
input   SRAM_WR, SRAM_RUN;
output  [31:0]  SRAM_RDATA;
output	UMORE, UMORE2LN;
output	DMA_IDLE;
/*output	UAD31O, UAD30O, UAD29O, UAD28O, UAD27O, UAD26O,
	UAD25O, UAD24O, UAD23O, UAD22O, UAD21O, UAD20O,
	UAD19O, UAD18O, UAD17O, UAD16O, UAD15O, UAD14O,
	UAD13O, UAD12O, UAD11O, UAD10O, UAD9O,  UAD8O,
	UAD7O,  UAD6O,  UAD5O,  UAD4O,  UAD3O,  UAD2O,
	UAD1O,  UAD0O;*/
output [31:0]   MA, MWD;

output	[31:0]	WPR;
output	MBE3_, MBE2_, MBE1_,MBE0_, CREQ, MRDY_, CACHEN,
	COMPL, MSWR, MRDMPLZ, XMITNULL,
	HCIGNT, TDMAEND, TXTHRESH;
/*input	PSADO31, PSADO30, PSADO29, PSADO28, PSADO27, PSADO26,
	PSADO25, PSADO24, PSADO23, PSADO22, PSADO21, PSADO20,
	PSADO19, PSADO18, PSADO17, PSADO16, PSADO15, PSADO14,
	PSADO13, PSADO12, PSADO11, PSADO10, PSADO9,  PSADO8,
	PSADO7,  PSADO6,  PSADO5,  PSADO4,  PSADO3,  PSADO2,
	PSADO1,  PSADO0;*/
input	AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I,
	AD23I, AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I,
	AD15I, AD14I, AD13I, AD12I, AD11I, AD10I, AD9I, AD8I,
	AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I;
input	[31:0]	BUFPTR1;
input	[19:0]	BUFPTR2;
input	[31:0]	HCIADR, HCIADD;
input	[10:0]	MAXLEN;
input	[7:0]	USBDAT;
output	[7:0]	HOSTDAT;
input	[7:0]	SLADDR;
input	CACHLN7, CACHLN6, CACHLN5, CACHLN4, CACHLN3, CACHLN2,
	CACHLN1, CACHLN0, CAHCFG_;
output	FEMPTY;
input	LATCHDAT, USBPOP;
input	QRXERR, MABORTS, TABORTR, BUSFREE, UGNTI_, //PMDSEL,
	MWRMEN, HCIREQ, HCICOMPL, HCIMWR, PMSTR, MADDR,
	PCI1WAIT, EOTQ, IN_DIR, RDYACK,
	/*UCBE3O_, UCBE2O_, UCBE1O_, UCBE0O_,*/ FCFG, HCIMRDY,
	/*TADOE, MADOE,*/ DIS_BURST, DISTXDLY2, BMUSM_RST_EN,
	DBUFERR, DISPFIFO, DISRXZERO, BUI_GO, DISPFIFO2,
	ENBMUSMRST, DISTXDLY, EOF,
	TEST_PACKET, SLAVEMODE, SLAVE_ACT, SLREAD, BIST_RUN,
	PCICLK, HRST_, BMUCRST_, CLK60M, HS_TRST_, ATPG_ENI;
output	/*UADOE_,*/ BOUNDRY;
output	[31:0]	MDO;
output	BIST_RUN_C, BIST_ERR_S, TESTPKTOK, DATARDY;

wire [31:0] FFRDPCI;
wire [3:0] FBE_;
wire [8:0] FCOUNT;

    zivc dnt08 ( .A(IN_DIR), .Y(TXFIFO) );
    zivc dnt09 ( .A(TXFIFO), .Y(RXFIFO) );
    zan2b DNTRXSTRT ( .A(LETSGO), .B(RXFIFO), .Y(RXSTRT) );
    zan2b DNTXMIT ( .A(LETSGO), .B(TXFIFO), .Y(XMITSTRT) );
    zckbufb dly6 ( .A(BUI_GO), .Y(BUISTRT) );
    zdl1b DD0 ( .A(MRDLY1), .Y(dd0) );
    zdl1b DD1 ( .A(BUISTRT), .Y(dd1) );
    zdffqb dly7 ( .D(dd1), .CK(PCICLK), .Q(MRDLY1) );
    zdffqb dly8 ( .D(dd0), .CK(PCICLK), .Q(LETSGO) );

    HS_BMUC HS_BMUC ( /*.UAD31O(UAD31O), .UAD30O(UAD30O), .UAD29O(UAD29O),
	.UAD28O(UAD28O), .UAD27O(UAD27O), .UAD26O(UAD26O), .UAD25O(UAD25O),
	.UAD24O(UAD24O), .UAD23O(UAD23O), .UAD22O(UAD22O), .UAD21O(UAD21O),
	.UAD20O(UAD20O), .UAD19O(UAD19O), .UAD18O(UAD18O), .UAD17O(UAD17O),
	.UAD16O(UAD16O), .UAD15O(UAD15O), .UAD14O(UAD14O), .UAD13O(UAD13O),
	.UAD12O(UAD12O), .UAD11O(UAD11O), .UAD10O(UAD10O), .UAD9O(UAD9O),
	.UAD8O(UAD8O), .UAD7O(UAD7O), .UAD6O(UAD6O), .UAD5O(UAD5O),
	.UAD4O(UAD4O), .UAD3O(UAD3O), .UAD2O(UAD2O), .UAD1O(UAD1O),
	.UAD0O(UAD0O),*/ .MA(MA), .MWD(MWD), .WPR(WPR), 
	.MBE3_(MBE3_), .MBE2_(MBE2_), .MBE1_(MBE1_), .MBE0_(MBE0_
	), .CREQ(CREQ), .MRDY_(MRDY_), .CACHEN(CACHEN), .COMPL(COMPL), .MSWR(
	MSWR), .MRDMPLZ(MRDMPLZ), .XMITNULL(XMITNULL), .PCIREAD(PCIREAD), 
	.PCIWRT(PCIWRT), .HCIGNT(HCIGNT), .RDMAEND(RDMAEND), .TDMAEND(TDMAEND)
	//, .TXTHRESH2(TXTHRESH2), .PSADO31(PSADO[31]), .PSADO30(PSADO[30]), 
	, .TXTHRESH(TXTHRESH), /*.PSADO31(PSADO31), .PSADO30(PSADO30), 
	.PSADO29(PSADO29), .PSADO28(PSADO28), .PSADO27(PSADO27), 
	.PSADO26(PSADO26), .PSADO25(PSADO25), .PSADO24(PSADO24), 
	.PSADO23(PSADO23), .PSADO22(PSADO22), .PSADO21(PSADO21), 
	.PSADO20(PSADO20), .PSADO19(PSADO19), .PSADO18(PSADO18), 
	.PSADO17(PSADO17), .PSADO16(PSADO16), .PSADO15(PSADO15), 
	.PSADO14(PSADO14), .PSADO13(PSADO13), .PSADO12(PSADO12), 
	.PSADO11(PSADO11), .PSADO10(PSADO10), .PSADO9(PSADO9), .PSADO8(
	PSADO8), .PSADO7(PSADO7), .PSADO6(PSADO6), .PSADO5(PSADO5), 
	.PSADO4(PSADO4), .PSADO3(PSADO3), .PSADO2(PSADO2), .PSADO1(
	PSADO1), .PSADO0(PSADO0),*/ .FFRDPCI(FFRDPCI),
	.BUFPTR1(BUFPTR1), .BUFPTR2({BUFPTR2, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
	1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
	.HCIADR(HCIADR), .HCIADD(HCIADD), .MAXLEN(MAXLEN),
	.CACHLN7(CACHLN7), .CACHLN6(CACHLN6), .CACHLN5(
	CACHLN5), .CACHLN4(CACHLN4), .CACHLN3(CACHLN3), .CACHLN2(
	CACHLN2), .CACHLN1(CACHLN1), .CACHLN0(CACHLN0), .CAHCFG_(CAHCFG_
	), .FBE_(FBE_),
	.RXPKTEND(RXPKTEND), .FEMPTY(FEMPTY), .FCOUNT(FCOUNT),
	.QRXERR(QRXERR), .MABORTS(MABORTS), .TABORTR(TABORTR), .XMITSTRT(
	XMITSTRT), .RXSTRT(RXSTRT), .BUSFREE(BUSFREE), .UGNTI_(UGNTI_), 
	/*.PMDSEL(PMDSEL),*/ .MWRMEN(MWRMEN), .HCIREQ(HCIREQ), .HCICOMPL(HCICOMPL)
	, .HCIMWR(HCIMWR), .PMSTR(PMSTR), .MADDR(MADDR), .PCI1WAIT(PCI1WAIT), 
	.EOTQ(EOTQ), .TXFIFO(TXFIFO), .RXFIFO(RXFIFO), .RDYACK(RDYACK), 
	/*.UCBE3O_(UCBE3O_), .UCBE2O_(UCBE2O_), .UCBE1O_(UCBE1O_), .UCBE0O_(
	UCBE0O_),*/ .FCFG(FCFG), .HCIMRDY(HCIMRDY), .PCICLK(PCICLK),
	.HRST_(BMUCRST_), .DISTXDLY(DISTXDLY),
	.EOF(EOF), .DISTXDLY2(DISTXDLY2), 
	.BMUSM_RST_EN(BMUSM_RST_EN), .DBUFERR(DBUFERR), .DISPFIFO(DISPFIFO), 
	.DISRXZERO(DISRXZERO), /*.ZEROLEN(ZEROLEN),*/ .BUI_GO(BUI_GO),
	.DISPFIFO2(DISPFIFO2), .ENBMUSMRST(ENBMUSMRST), .TADOE(1'b1),
	/*.MADOE(1'b1), .UADOE_(UADOE_),*/ .BOUNDRY(BOUNDRY),
	.DIS_BURST(DIS_BURST), .DMA_IDLE(DMA_IDLE),
	.UMORE(UMORE), .UMORE2LN(UMORE2LN), .ATPG_ENI(ATPG_ENI),
	.FIFO_OK(FIFO_OK) );

    HS_PER_FIFO HS_FIFO ( .FFRDPCI(FFRDPCI), .HOSTDAT(HOSTDAT),
	.FCOUNT(FCOUNT), .FFULL(FFULL), .FEMPTY(FEMPTY), .FBE_(FBE_),
	.RXPKTEND(RXPKTEND), .USBDAT(USBDAT), .ADI({AD31I,
        AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I, AD23I, AD22I, AD21I,
        AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, AD14I, AD13I, AD12I, AD11I,
        AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I}),
	.BUISTRT(BUISTRT), .XMITSTRT(XMITSTRT), .RXFIFO(RXFIFO),
	.LATCHDAT(LATCHDAT), .USBPOP(USBPOP), .PCIWRT(PCIWRT), 
	.PCIREAD(PCIREAD), .EOTQ(EOTQ), .RDMAEND(RDMAEND), .WPR1(WPR[1]),
	.WPR0(WPR[0]), //.UCBEO_({UCBE3O_, UCBE2O_, UCBE1O_, UCBE0O_}),
	.UCBEO_({MBE3_, MBE2_, MBE1_, MBE0_}),
	.PCICLK(PCICLK), .CLK60M(CLK60M), .HRST_(HRST_), .TRST_(HS_TRST_),
	.RXSTRT(RXSTRT), .FIFO_OK(FIFO_OK), .TDMAEND(TDMAEND),
	.RXERR(QRXERR), .TEST_PACKET(TEST_PACKET), .TESTPKTOK(TESTPKTOK),
	.SLAVEMODE(SLAVEMODE), .SLADDR(SLADDR), .DATARDY(DATARDY),
	.SLREAD(SLREAD), .MDO(MDO), .SLAVE_ACT(SLAVE_ACT),
	.BIST_RUN(BIST_RUN), .BIST_RUN_C(BIST_RUN_C),
        .BIST_ERR_S(BIST_ERR_S), .ATPG_ENI(ATPG_ENI),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_ID(SRAM_ID), .SRAM_WR(SRAM_WR),
        .SRAM_RUN(SRAM_RUN), .SRAM_RDATA(SRAM_RDATA),
	.ATPG_CLK(ATPG_CLK) );

endmodule

// USB 2.0 HS asynchronous DMA controller
module HS_ASYNC_DMA ( /*UAD31O, UAD30O, UAD29O, UAD28O, UAD27O, UAD26O,
		UAD25O, UAD24O, UAD23O, UAD22O, UAD21O, UAD20O,
                UAD19O, UAD18O, UAD17O, UAD16O, UAD15O, UAD14O,
                UAD13O, UAD12O, UAD11O, UAD10O, UAD9O,  UAD8O,
                UAD7O,  UAD6O,  UAD5O,  UAD4O,  UAD3O,  UAD2O,
                UAD1O,  UAD0O,*/
		MA, MWD, WPR,
		MBE3_, MBE2_, MBE1_,MBE0_, CREQ, MRDY_, CACHEN,
		COMPL, MSWR, MRDMPLZ, XMITNULL,
		UMORE, UMORE2LN,
                HCIGNT, TDMAEND, TXTHRESH,
		/*PSADO31, PSADO30, PSADO29, PSADO28, PSADO27, PSADO26,
                PSADO25, PSADO24, PSADO23, PSADO22, PSADO21, PSADO20,
                PSADO19, PSADO18, PSADO17, PSADO16, PSADO15, PSADO14,
                PSADO13, PSADO12, PSADO11, PSADO10, PSADO9,  PSADO8,
                PSADO7,  PSADO6,  PSADO5,  PSADO4,  PSADO3,  PSADO2,
                PSADO1,  PSADO0,*/
		AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I,
		AD23I, AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I,
		AD15I, AD14I, AD13I, AD12I, AD11I, AD10I, AD9I, AD8I,
		AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I,
		BUFPTR1, BUFPTR2, HCIADR, HCIADD, MAXLEN,
		USBDAT, LATCHDAT, USBPOP, HOSTDAT,
		CACHLN7,  CACHLN6,  CACHLN5,  CACHLN4,  CACHLN3,  CACHLN2,
                CACHLN1,  CACHLN0, CAHCFG_,
		FEMPTY,
		QRXERR, MABORTS, TABORTR,
		BUSFREE , UGNTI_, /*PMDSEL,*/ MWRMEN,
		HCIREQ, HCICOMPL, HCIMWR, PMSTR, MADDR, PCI1WAIT,
		EOTQ, IN_DIR, RDYACK,
		//UCBE3O_, UCBE2O_, UCBE1O_,UCBE0O_,
		FCFG, HCIMRDY,
		DISTXDLY, EOF,
		DISTXDLY2, BMUSM_RST_EN, DBUFERR, DISPFIFO,
		DISRXZERO, BUI_GO, DISPFIFO2,
		ENBMUSMRST, /*TADOE, MADOE, UADOE_,*/ BOUNDRY, DIS_BURST,
		TEST_PACKET, SLAVEMODE, SLAVE_ACT, SLADDR, SLREAD,
		BIST_RUN, BIST_RUN_C, BIST_ERR_S, TESTPKTOK, DATARDY,
		MDO, PCICLK, HRST_, BMUCRST_, CLK60M, HS_TRST_, DMA_IDLE,
		ATPG_ENI, BIST_PATTERN, SRAM_ADDR, SRAM_SEL, SRAM_WR, SRAM_RUN,
                SRAM_ID, SRAM_RDATA, ATPG_CLK
		);
input	ATPG_CLK;
input   [31:0]  BIST_PATTERN;
input   [8:0]   SRAM_ADDR;
input   [1:0]   SRAM_SEL, SRAM_ID;
input   SRAM_WR, SRAM_RUN;
output  [31:0]  SRAM_RDATA;
output	UMORE, UMORE2LN;
output	DMA_IDLE;
/*output	UAD31O, UAD30O, UAD29O, UAD28O, UAD27O, UAD26O,
	UAD25O, UAD24O, UAD23O, UAD22O, UAD21O, UAD20O,
	UAD19O, UAD18O, UAD17O, UAD16O, UAD15O, UAD14O,
	UAD13O, UAD12O, UAD11O, UAD10O, UAD9O,  UAD8O,
	UAD7O,  UAD6O,  UAD5O,  UAD4O,  UAD3O,  UAD2O,
	UAD1O,  UAD0O;*/
output [31:0]   MA, MWD;

output	[31:0]	WPR;
output	MBE3_, MBE2_, MBE1_,MBE0_, CREQ, MRDY_, CACHEN,
	COMPL, MSWR, MRDMPLZ, XMITNULL,
	HCIGNT, TDMAEND, TXTHRESH;
/*input	PSADO31, PSADO30, PSADO29, PSADO28, PSADO27, PSADO26,
	PSADO25, PSADO24, PSADO23, PSADO22, PSADO21, PSADO20,
	PSADO19, PSADO18, PSADO17, PSADO16, PSADO15, PSADO14,
	PSADO13, PSADO12, PSADO11, PSADO10, PSADO9,  PSADO8,
	PSADO7,  PSADO6,  PSADO5,  PSADO4,  PSADO3,  PSADO2,
	PSADO1,  PSADO0;*/
input	AD31I, AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I,
	AD23I, AD22I, AD21I, AD20I, AD19I, AD18I, AD17I, AD16I,
	AD15I, AD14I, AD13I, AD12I, AD11I, AD10I, AD9I, AD8I,
	AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I;
input	[31:0]	BUFPTR1;
input	[19:0]	BUFPTR2;
input	[31:0]	HCIADR, HCIADD;
input	[10:0]	MAXLEN;
input	[7:0]	USBDAT;
output	[7:0]	HOSTDAT;
input	[7:0]	SLADDR;
input	CACHLN7, CACHLN6, CACHLN5, CACHLN4, CACHLN3, CACHLN2,
	CACHLN1, CACHLN0, CAHCFG_;
output	FEMPTY;
input	LATCHDAT, USBPOP;
input	QRXERR, MABORTS, TABORTR, BUSFREE, UGNTI_, //PMDSEL,
	MWRMEN, HCIREQ, HCICOMPL, HCIMWR, PMSTR, MADDR,
	PCI1WAIT, EOTQ, IN_DIR, RDYACK,
	/*UCBE3O_, UCBE2O_, UCBE1O_, UCBE0O_,*/ FCFG, HCIMRDY,
	/*TADOE, MADOE,*/ DIS_BURST, DISTXDLY2, BMUSM_RST_EN,
	DBUFERR, DISPFIFO, DISRXZERO, BUI_GO, DISPFIFO2,
	ENBMUSMRST, DISTXDLY, EOF,
	TEST_PACKET, SLAVEMODE, SLAVE_ACT, SLREAD, BIST_RUN,
	PCICLK, HRST_, BMUCRST_, CLK60M, HS_TRST_, ATPG_ENI;
output	/*UADOE_,*/ BOUNDRY;
output	[31:0]	MDO;
output	BIST_RUN_C, BIST_ERR_S, TESTPKTOK, DATARDY;

wire [31:0] FFRDPCI;
wire [3:0] FBE_;
wire [8:0] FCOUNT;

    zivc dnt08 ( .A(IN_DIR), .Y(TXFIFO) );
    zivc dnt09 ( .A(TXFIFO), .Y(RXFIFO) );
    zan2b DNTRXSTRT ( .A(LETSGO), .B(RXFIFO), .Y(RXSTRT) );
    zan2b DNTXMIT ( .A(LETSGO), .B(TXFIFO), .Y(XMITSTRT) );
    zckbufb dly6 ( .A(BUI_GO), .Y(BUISTRT) );
    zdl1b DD0 ( .A(MRDLY1), .Y(dd0) );
    zdl1b DD1 ( .A(BUISTRT), .Y(dd1) );
    zdffqb dly7 ( .D(dd1), .CK(PCICLK), .Q(MRDLY1) );
    zdffqb dly8 ( .D(dd0), .CK(PCICLK), .Q(LETSGO) );

    HS_BMUC HS_BMUC ( /*.UAD31O(UAD31O), .UAD30O(UAD30O), .UAD29O(UAD29O),
	.UAD28O(UAD28O), .UAD27O(UAD27O), .UAD26O(UAD26O), .UAD25O(UAD25O),
	.UAD24O(UAD24O), .UAD23O(UAD23O), .UAD22O(UAD22O), .UAD21O(UAD21O),
	.UAD20O(UAD20O), .UAD19O(UAD19O), .UAD18O(UAD18O), .UAD17O(UAD17O),
	.UAD16O(UAD16O), .UAD15O(UAD15O), .UAD14O(UAD14O), .UAD13O(UAD13O),
	.UAD12O(UAD12O), .UAD11O(UAD11O), .UAD10O(UAD10O), .UAD9O(UAD9O),
	.UAD8O(UAD8O), .UAD7O(UAD7O), .UAD6O(UAD6O), .UAD5O(UAD5O),
	.UAD4O(UAD4O), .UAD3O(UAD3O), .UAD2O(UAD2O), .UAD1O(UAD1O),
	.UAD0O(UAD0O),*/ .MA(MA), .MWD(MWD), .WPR(WPR), 
	.MBE3_(MBE3_), .MBE2_(MBE2_), .MBE1_(MBE1_), .MBE0_(MBE0_
	), .CREQ(CREQ), .MRDY_(MRDY_), .CACHEN(CACHEN), .COMPL(COMPL), .MSWR(
	MSWR), .MRDMPLZ(MRDMPLZ), .XMITNULL(XMITNULL), .PCIREAD(PCIREAD), 
	.PCIWRT(PCIWRT), .HCIGNT(HCIGNT), .RDMAEND(RDMAEND), .TDMAEND(TDMAEND)
	//, .TXTHRESH2(TXTHRESH2), .PSADO31(PSADO[31]), .PSADO30(PSADO[30]), 
	, .TXTHRESH(TXTHRESH), /*.PSADO31(PSADO31), .PSADO30(PSADO30), 
	.PSADO29(PSADO29), .PSADO28(PSADO28), .PSADO27(PSADO27), 
	.PSADO26(PSADO26), .PSADO25(PSADO25), .PSADO24(PSADO24), 
	.PSADO23(PSADO23), .PSADO22(PSADO22), .PSADO21(PSADO21), 
	.PSADO20(PSADO20), .PSADO19(PSADO19), .PSADO18(PSADO18), 
	.PSADO17(PSADO17), .PSADO16(PSADO16), .PSADO15(PSADO15), 
	.PSADO14(PSADO14), .PSADO13(PSADO13), .PSADO12(PSADO12), 
	.PSADO11(PSADO11), .PSADO10(PSADO10), .PSADO9(PSADO9), .PSADO8(
	PSADO8), .PSADO7(PSADO7), .PSADO6(PSADO6), .PSADO5(PSADO5), 
	.PSADO4(PSADO4), .PSADO3(PSADO3), .PSADO2(PSADO2), .PSADO1(
	PSADO1), .PSADO0(PSADO0),*/ .FFRDPCI(FFRDPCI),
	.BUFPTR1(BUFPTR1), .BUFPTR2({BUFPTR2, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
	1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
	.HCIADR(HCIADR), .HCIADD(HCIADD), .MAXLEN(MAXLEN),
	.CACHLN7(CACHLN7), .CACHLN6(CACHLN6), .CACHLN5(
	CACHLN5), .CACHLN4(CACHLN4), .CACHLN3(CACHLN3), .CACHLN2(
	CACHLN2), .CACHLN1(CACHLN1), .CACHLN0(CACHLN0), .CAHCFG_(CAHCFG_
	), .FBE_(FBE_),
	.RXPKTEND(RXPKTEND), .FEMPTY(FEMPTY), .FCOUNT(FCOUNT),
	.QRXERR(QRXERR), .MABORTS(MABORTS), .TABORTR(TABORTR), .XMITSTRT(
	XMITSTRT), .RXSTRT(RXSTRT), .BUSFREE(BUSFREE), .UGNTI_(UGNTI_), 
	/*.PMDSEL(PMDSEL),*/ .MWRMEN(MWRMEN), .HCIREQ(HCIREQ), .HCICOMPL(HCICOMPL)
	, .HCIMWR(HCIMWR), .PMSTR(PMSTR), .MADDR(MADDR), .PCI1WAIT(PCI1WAIT), 
	.EOTQ(EOTQ), .TXFIFO(TXFIFO), .RXFIFO(RXFIFO), .RDYACK(RDYACK), 
	/*.UCBE3O_(UCBE3O_), .UCBE2O_(UCBE2O_), .UCBE1O_(UCBE1O_), .UCBE0O_(
	UCBE0O_),*/ .FCFG(FCFG), .HCIMRDY(HCIMRDY), .PCICLK(PCICLK),
	.HRST_(BMUCRST_), .DISTXDLY(DISTXDLY),
	.EOF(EOF), .DISTXDLY2(DISTXDLY2), 
	.BMUSM_RST_EN(BMUSM_RST_EN), .DBUFERR(DBUFERR), .DISPFIFO(DISPFIFO), 
	.DISRXZERO(DISRXZERO), /*.ZEROLEN(ZEROLEN),*/ .BUI_GO(BUI_GO),
	.DISPFIFO2(DISPFIFO2), .ENBMUSMRST(ENBMUSMRST), .TADOE(1'b1),
	/*.MADOE(1'b1), .UADOE_(UADOE_),*/ .BOUNDRY(BOUNDRY),
	.DIS_BURST(DIS_BURST), .DMA_IDLE(DMA_IDLE),
	.UMORE(UMORE), .UMORE2LN(UMORE2LN), .ATPG_ENI(ATPG_ENI),
	.FIFO_OK(FIFO_OK) );

    HS_ASYNC_FIFO HS_FIFO ( .FFRDPCI(FFRDPCI), .HOSTDAT(HOSTDAT),
	.FCOUNT(FCOUNT), .FFULL(FFULL), .FEMPTY(FEMPTY), .FBE_(FBE_),
	.RXPKTEND(RXPKTEND), .USBDAT(USBDAT), .ADI({AD31I,
        AD30I, AD29I, AD28I, AD27I, AD26I, AD25I, AD24I, AD23I, AD22I, AD21I,
        AD20I, AD19I, AD18I, AD17I, AD16I, AD15I, AD14I, AD13I, AD12I, AD11I,
        AD10I, AD9I, AD8I, AD7I, AD6I, AD5I, AD4I, AD3I, AD2I, AD1I, AD0I}),
	.BUISTRT(BUISTRT), .XMITSTRT(XMITSTRT), .RXFIFO(RXFIFO),
	.LATCHDAT(LATCHDAT), .USBPOP(USBPOP), .PCIWRT(PCIWRT), 
	.PCIREAD(PCIREAD), .EOTQ(EOTQ), .RDMAEND(RDMAEND), .WPR1(WPR[1]),
	.WPR0(WPR[0]), //.UCBEO_({UCBE3O_, UCBE2O_, UCBE1O_, UCBE0O_}),
	.UCBEO_({MBE3_, MBE2_, MBE1_, MBE0_}),
	.PCICLK(PCICLK), .CLK60M(CLK60M), .HRST_(HRST_), .TRST_(HS_TRST_),
	.RXSTRT(RXSTRT), .FIFO_OK(FIFO_OK), .TDMAEND(TDMAEND),
	.RXERR(QRXERR), .TEST_PACKET(TEST_PACKET), .TESTPKTOK(TESTPKTOK),
	.SLAVEMODE(SLAVEMODE), .SLADDR(SLADDR), .DATARDY(DATARDY),
	.SLREAD(SLREAD), .MDO(MDO), .SLAVE_ACT(SLAVE_ACT),
	.BIST_RUN(BIST_RUN), .BIST_RUN_C(BIST_RUN_C),
        .BIST_ERR_S(BIST_ERR_S), .ATPG_ENI(ATPG_ENI),
	.BIST_PATTERN(BIST_PATTERN), .SRAM_ADDR(SRAM_ADDR),
        .SRAM_SEL(SRAM_SEL), .SRAM_ID(SRAM_ID), .SRAM_WR(SRAM_WR),
        .SRAM_RUN(SRAM_RUN), .SRAM_RDATA(SRAM_RDATA),
	.ATPG_CLK(ATPG_CLK) );

endmodule

